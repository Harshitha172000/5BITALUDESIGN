magic
tech scmos
timestamp 1606902023
<< rotate >>
rect 155 223 166 225
rect 432 223 443 225
rect 708 223 719 225
rect 985 223 996 225
rect 132 219 134 221
rect 155 216 169 223
rect 409 219 411 221
rect 432 216 446 223
rect 685 219 687 221
rect 708 216 722 223
rect 962 219 964 221
rect 985 216 999 223
rect 158 214 169 216
rect 435 214 446 216
rect 711 214 722 216
rect 988 214 999 216
rect 155 79 166 81
rect 432 79 443 81
rect 708 79 719 81
rect 985 79 996 81
rect 132 75 134 77
rect 155 72 169 79
rect 409 75 411 77
rect 432 72 446 79
rect 685 75 687 77
rect 708 72 722 79
rect 962 75 964 77
rect 985 72 999 79
rect 158 70 169 72
rect 435 70 446 72
rect 711 70 722 72
rect 988 70 999 72
<< ab >>
rect -290 288 -289 360
rect -285 0 -221 360
rect -217 346 -40 360
rect -217 342 -215 346
rect -213 342 -43 346
rect -41 342 -40 346
rect -217 234 -40 342
rect -217 230 -215 234
rect -213 230 -43 234
rect -41 230 -40 234
rect -217 202 -40 230
rect -217 198 -215 202
rect -213 198 -43 202
rect -41 198 -40 202
rect -217 90 -40 198
rect -217 86 -215 90
rect -213 86 -43 90
rect -41 86 -40 90
rect -217 58 -40 86
rect -217 54 -215 58
rect -213 54 -43 58
rect -41 54 -40 58
rect -217 0 -40 54
rect -38 1 3 360
rect -39 0 3 1
rect 5 346 262 360
rect 5 342 87 346
rect 89 342 259 346
rect 261 342 262 346
rect 5 234 262 342
rect 5 230 87 234
rect 89 230 259 234
rect 261 230 262 234
rect 5 202 262 230
rect 5 198 87 202
rect 89 198 259 202
rect 261 198 262 202
rect 5 90 262 198
rect 5 86 87 90
rect 89 86 259 90
rect 261 86 262 90
rect 5 58 262 86
rect 5 54 87 58
rect 89 54 259 58
rect 261 54 262 58
rect 5 0 262 54
rect 264 249 305 360
rect 264 246 306 249
rect 264 105 305 246
rect 264 102 306 105
rect 264 0 305 102
rect 312 0 352 360
rect 361 346 539 360
rect 361 342 364 346
rect 366 342 536 346
rect 538 342 539 346
rect 361 234 539 342
rect 361 230 364 234
rect 366 230 536 234
rect 538 230 539 234
rect 361 202 539 230
rect 361 198 364 202
rect 366 198 536 202
rect 538 198 539 202
rect 361 90 539 198
rect 361 86 364 90
rect 366 86 536 90
rect 538 86 539 90
rect 361 58 539 86
rect 361 54 364 58
rect 366 54 536 58
rect 538 54 539 58
rect 361 0 539 54
rect 541 249 582 360
rect 541 246 583 249
rect 541 105 582 246
rect 541 102 583 105
rect 541 0 582 102
rect 589 1 629 360
rect 637 346 815 360
rect 637 342 640 346
rect 642 342 812 346
rect 814 342 815 346
rect 637 234 815 342
rect 637 230 640 234
rect 642 230 812 234
rect 814 230 815 234
rect 637 202 815 230
rect 637 198 640 202
rect 642 198 812 202
rect 814 198 815 202
rect 637 90 815 198
rect 637 86 640 90
rect 642 86 812 90
rect 814 86 815 90
rect 637 58 815 86
rect 637 54 640 58
rect 642 54 812 58
rect 814 54 815 58
rect 637 1 815 54
rect 817 249 858 360
rect 817 246 859 249
rect 817 105 858 246
rect 817 102 859 105
rect 817 1 858 102
rect 865 1 905 360
rect 914 346 1092 360
rect 914 342 917 346
rect 919 342 1089 346
rect 1091 342 1092 346
rect 914 234 1092 342
rect 914 230 917 234
rect 919 230 1089 234
rect 1091 230 1092 234
rect 914 202 1092 230
rect 914 198 917 202
rect 919 198 1089 202
rect 1091 198 1092 202
rect 914 90 1092 198
rect 914 86 917 90
rect 919 86 1089 90
rect 1091 86 1092 90
rect 914 58 1092 86
rect 914 54 917 58
rect 919 54 1089 58
rect 1091 54 1092 58
rect 914 1 1092 54
rect 1094 249 1135 360
rect 1094 246 1136 249
rect 1094 105 1135 246
rect 1094 102 1136 105
rect 1094 1 1135 102
rect 589 0 1135 1
rect -158 -71 154 0
rect 160 -71 225 0
rect 226 -71 247 0
rect 248 -71 289 0
rect 291 -71 553 0
rect 555 -71 597 0
rect 599 -71 1071 0
rect 1075 -71 1131 0
<< nwell >>
rect -290 364 201 365
rect 250 364 478 365
rect 527 364 754 365
rect 803 364 1031 365
rect 1080 364 1136 365
rect -290 320 1136 364
rect -290 176 1136 256
rect -290 32 1136 112
rect -158 -76 1136 -31
<< pwell >>
rect -290 256 1136 320
rect -290 112 1136 176
rect -290 -5 1136 32
rect -181 -7 1136 -5
rect -158 -31 1136 -7
<< poly >>
rect -268 354 -266 358
rect -283 329 -277 331
rect -283 327 -281 329
rect -279 327 -277 329
rect -232 354 -230 358
rect -208 354 -206 358
rect -252 345 -250 349
rect -242 345 -240 349
rect -185 351 -183 356
rect -178 351 -176 356
rect -160 354 -158 358
rect -150 354 -148 358
rect -140 354 -138 358
rect -118 354 -116 358
rect -108 354 -106 358
rect -98 354 -96 358
rect -195 342 -193 347
rect -283 325 -277 327
rect -279 324 -277 325
rect -268 324 -266 327
rect -252 324 -250 327
rect -279 322 -266 324
rect -260 322 -250 324
rect -242 323 -240 327
rect -232 324 -230 327
rect -276 314 -274 322
rect -260 318 -258 322
rect -267 316 -258 318
rect -246 321 -240 323
rect -246 319 -244 321
rect -242 319 -240 321
rect -246 317 -240 319
rect -236 322 -230 324
rect -236 320 -234 322
rect -232 320 -230 322
rect -236 318 -230 320
rect -267 314 -265 316
rect -263 314 -258 316
rect -267 312 -258 314
rect -242 314 -240 317
rect -260 309 -258 312
rect -250 309 -248 313
rect -242 312 -238 314
rect -240 309 -238 312
rect -233 309 -231 318
rect -208 316 -206 329
rect -195 326 -193 329
rect -80 351 -78 356
rect -73 351 -71 356
rect -50 354 -48 358
rect -29 354 -27 358
rect -22 354 -20 358
rect -63 342 -61 347
rect -9 344 -7 349
rect 14 347 16 352
rect 24 347 26 352
rect 94 354 96 358
rect -29 330 -27 333
rect -63 326 -61 329
rect -202 324 -193 326
rect -202 322 -200 324
rect -198 322 -196 324
rect -185 323 -183 326
rect -178 323 -176 326
rect -160 323 -158 326
rect -150 323 -148 326
rect -140 323 -138 326
rect -118 323 -116 326
rect -108 323 -106 326
rect -98 323 -96 326
rect -80 323 -78 326
rect -73 323 -71 326
rect -63 324 -54 326
rect -202 320 -196 322
rect -208 314 -202 316
rect -208 312 -206 314
rect -204 312 -202 314
rect -208 310 -202 312
rect -276 302 -274 305
rect -276 300 -271 302
rect -273 292 -271 300
rect -260 296 -258 300
rect -250 292 -248 300
rect -208 307 -206 310
rect -198 307 -196 320
rect -188 321 -182 323
rect -188 319 -186 321
rect -184 319 -182 321
rect -188 317 -182 319
rect -178 321 -156 323
rect -178 319 -167 321
rect -165 319 -160 321
rect -158 319 -156 321
rect -178 317 -156 319
rect -152 321 -146 323
rect -152 319 -150 321
rect -148 319 -146 321
rect -152 317 -146 319
rect -142 321 -136 323
rect -142 319 -140 321
rect -138 319 -136 321
rect -142 317 -136 319
rect -120 321 -114 323
rect -120 319 -118 321
rect -116 319 -114 321
rect -120 317 -114 319
rect -110 321 -104 323
rect -110 319 -108 321
rect -106 319 -104 321
rect -110 317 -104 319
rect -100 321 -78 323
rect -100 319 -98 321
rect -96 319 -91 321
rect -89 319 -78 321
rect -100 317 -78 319
rect -74 321 -68 323
rect -74 319 -72 321
rect -70 319 -68 321
rect -74 317 -68 319
rect -188 314 -186 317
rect -178 314 -176 317
rect -158 314 -156 317
rect -151 314 -149 317
rect -240 292 -238 297
rect -233 292 -231 297
rect -273 290 -248 292
rect -208 290 -206 294
rect -198 292 -196 297
rect -188 295 -186 300
rect -178 295 -176 300
rect -140 308 -138 317
rect -118 308 -116 317
rect -107 314 -105 317
rect -100 314 -98 317
rect -80 314 -78 317
rect -70 314 -68 317
rect -60 322 -58 324
rect -56 322 -54 324
rect -60 320 -54 322
rect -60 307 -58 320
rect -50 316 -48 329
rect -33 328 -27 330
rect -33 326 -31 328
rect -29 326 -27 328
rect -33 324 -27 326
rect -54 314 -48 316
rect -29 314 -27 324
rect -22 323 -20 333
rect 34 345 36 349
rect 54 347 56 352
rect 64 347 66 352
rect 14 331 16 334
rect 10 329 16 331
rect 10 327 12 329
rect 14 327 16 329
rect -9 323 -7 326
rect 10 325 16 327
rect -23 321 -17 323
rect -23 319 -21 321
rect -19 319 -17 321
rect -23 317 -17 319
rect -13 321 -7 323
rect -13 319 -11 321
rect -9 319 -7 321
rect -13 317 -7 319
rect -19 314 -17 317
rect -9 314 -7 317
rect -54 312 -52 314
rect -50 312 -48 314
rect -54 310 -48 312
rect -50 307 -48 310
rect -80 295 -78 300
rect -70 295 -68 300
rect -158 290 -156 294
rect -151 290 -149 294
rect -140 290 -138 294
rect -118 290 -116 294
rect -107 290 -105 294
rect -100 290 -98 294
rect -60 292 -58 297
rect -29 303 -27 308
rect -19 303 -17 308
rect 14 312 16 325
rect 24 323 26 334
rect 74 345 76 349
rect 54 331 56 334
rect 50 329 56 331
rect 50 327 52 329
rect 54 327 56 329
rect 34 323 36 327
rect 50 325 56 327
rect 20 321 26 323
rect 20 319 22 321
rect 24 319 26 321
rect 20 317 26 319
rect 30 321 36 323
rect 30 319 32 321
rect 34 319 36 321
rect 30 317 36 319
rect 21 312 23 317
rect 34 312 36 317
rect 54 312 56 325
rect 64 323 66 334
rect 117 351 119 356
rect 124 351 126 356
rect 142 354 144 358
rect 152 354 154 358
rect 162 354 164 358
rect 184 354 186 358
rect 194 354 196 358
rect 204 354 206 358
rect 107 342 109 347
rect 74 323 76 327
rect 60 321 66 323
rect 60 319 62 321
rect 64 319 66 321
rect 60 317 66 319
rect 70 321 76 323
rect 70 319 72 321
rect 74 319 76 321
rect 70 317 76 319
rect 61 312 63 317
rect 74 312 76 317
rect 94 316 96 329
rect 107 326 109 329
rect 222 351 224 356
rect 229 351 231 356
rect 252 354 254 358
rect 273 354 275 358
rect 280 354 282 358
rect 239 342 241 347
rect 371 354 373 358
rect 293 344 295 349
rect 321 347 323 352
rect 331 347 333 352
rect 273 330 275 333
rect 239 326 241 329
rect 100 324 109 326
rect 100 322 102 324
rect 104 322 106 324
rect 117 323 119 326
rect 124 323 126 326
rect 142 323 144 326
rect 152 323 154 326
rect 162 323 164 326
rect 184 323 186 326
rect 194 323 196 326
rect 204 323 206 326
rect 222 323 224 326
rect 229 323 231 326
rect 239 324 248 326
rect 100 320 106 322
rect 94 314 100 316
rect 94 312 96 314
rect 98 312 100 314
rect -9 300 -7 305
rect 14 296 16 301
rect 21 296 23 301
rect -50 290 -48 294
rect 34 299 36 303
rect 94 310 100 312
rect 94 307 96 310
rect 104 307 106 320
rect 114 321 120 323
rect 114 319 116 321
rect 118 319 120 321
rect 114 317 120 319
rect 124 321 146 323
rect 124 319 135 321
rect 137 319 142 321
rect 144 319 146 321
rect 124 317 146 319
rect 150 321 156 323
rect 150 319 152 321
rect 154 319 156 321
rect 150 317 156 319
rect 160 321 166 323
rect 160 319 162 321
rect 164 319 166 321
rect 160 317 166 319
rect 182 321 188 323
rect 182 319 184 321
rect 186 319 188 321
rect 182 317 188 319
rect 192 321 198 323
rect 192 319 194 321
rect 196 319 198 321
rect 192 317 198 319
rect 202 321 224 323
rect 202 319 204 321
rect 206 319 211 321
rect 213 319 224 321
rect 202 317 224 319
rect 228 321 234 323
rect 228 319 230 321
rect 232 319 234 321
rect 228 317 234 319
rect 114 314 116 317
rect 124 314 126 317
rect 144 314 146 317
rect 151 314 153 317
rect 54 296 56 301
rect 61 296 63 301
rect 74 299 76 303
rect 94 290 96 294
rect 104 292 106 297
rect 114 295 116 300
rect 124 295 126 300
rect 162 308 164 317
rect 184 308 186 317
rect 195 314 197 317
rect 202 314 204 317
rect 222 314 224 317
rect 232 314 234 317
rect 242 322 244 324
rect 246 322 248 324
rect 242 320 248 322
rect 242 307 244 320
rect 252 316 254 329
rect 269 328 275 330
rect 269 326 271 328
rect 273 326 275 328
rect 269 324 275 326
rect 248 314 254 316
rect 273 314 275 324
rect 280 323 282 333
rect 341 345 343 349
rect 321 331 323 334
rect 317 329 323 331
rect 317 327 319 329
rect 321 327 323 329
rect 293 323 295 326
rect 317 325 323 327
rect 279 321 285 323
rect 279 319 281 321
rect 283 319 285 321
rect 279 317 285 319
rect 289 321 295 323
rect 289 319 291 321
rect 293 319 295 321
rect 289 317 295 319
rect 283 314 285 317
rect 293 314 295 317
rect 248 312 250 314
rect 252 312 254 314
rect 248 310 254 312
rect 252 307 254 310
rect 222 295 224 300
rect 232 295 234 300
rect 144 290 146 294
rect 151 290 153 294
rect 162 290 164 294
rect 184 290 186 294
rect 195 290 197 294
rect 202 290 204 294
rect 242 292 244 297
rect 273 303 275 308
rect 283 303 285 308
rect 321 312 323 325
rect 331 323 333 334
rect 394 351 396 356
rect 401 351 403 356
rect 419 354 421 358
rect 429 354 431 358
rect 439 354 441 358
rect 461 354 463 358
rect 471 354 473 358
rect 481 354 483 358
rect 384 342 386 347
rect 341 323 343 327
rect 327 321 333 323
rect 327 319 329 321
rect 331 319 333 321
rect 327 317 333 319
rect 337 321 343 323
rect 337 319 339 321
rect 341 319 343 321
rect 337 317 343 319
rect 328 312 330 317
rect 341 312 343 317
rect 371 316 373 329
rect 384 326 386 329
rect 499 351 501 356
rect 506 351 508 356
rect 529 354 531 358
rect 550 354 552 358
rect 557 354 559 358
rect 516 342 518 347
rect 647 354 649 358
rect 570 344 572 349
rect 598 347 600 352
rect 608 347 610 352
rect 550 330 552 333
rect 516 326 518 329
rect 377 324 386 326
rect 377 322 379 324
rect 381 322 383 324
rect 394 323 396 326
rect 401 323 403 326
rect 419 323 421 326
rect 429 323 431 326
rect 439 323 441 326
rect 461 323 463 326
rect 471 323 473 326
rect 481 323 483 326
rect 499 323 501 326
rect 506 323 508 326
rect 516 324 525 326
rect 377 320 383 322
rect 371 314 377 316
rect 371 312 373 314
rect 375 312 377 314
rect 293 300 295 305
rect 371 310 377 312
rect 371 307 373 310
rect 381 307 383 320
rect 391 321 397 323
rect 391 319 393 321
rect 395 319 397 321
rect 391 317 397 319
rect 401 321 423 323
rect 401 319 412 321
rect 414 319 419 321
rect 421 319 423 321
rect 401 317 423 319
rect 427 321 433 323
rect 427 319 429 321
rect 431 319 433 321
rect 427 317 433 319
rect 437 321 443 323
rect 437 319 439 321
rect 441 319 443 321
rect 437 317 443 319
rect 459 321 465 323
rect 459 319 461 321
rect 463 319 465 321
rect 459 317 465 319
rect 469 321 475 323
rect 469 319 471 321
rect 473 319 475 321
rect 469 317 475 319
rect 479 321 501 323
rect 479 319 481 321
rect 483 319 488 321
rect 490 319 501 321
rect 479 317 501 319
rect 505 321 511 323
rect 505 319 507 321
rect 509 319 511 321
rect 505 317 511 319
rect 391 314 393 317
rect 401 314 403 317
rect 421 314 423 317
rect 428 314 430 317
rect 321 296 323 301
rect 328 296 330 301
rect 252 290 254 294
rect 341 299 343 303
rect 371 290 373 294
rect 381 292 383 297
rect 391 295 393 300
rect 401 295 403 300
rect 439 308 441 317
rect 461 308 463 317
rect 472 314 474 317
rect 479 314 481 317
rect 499 314 501 317
rect 509 314 511 317
rect 519 322 521 324
rect 523 322 525 324
rect 519 320 525 322
rect 519 307 521 320
rect 529 316 531 329
rect 546 328 552 330
rect 546 326 548 328
rect 550 326 552 328
rect 546 324 552 326
rect 525 314 531 316
rect 550 314 552 324
rect 557 323 559 333
rect 618 345 620 349
rect 598 331 600 334
rect 594 329 600 331
rect 594 327 596 329
rect 598 327 600 329
rect 570 323 572 326
rect 594 325 600 327
rect 556 321 562 323
rect 556 319 558 321
rect 560 319 562 321
rect 556 317 562 319
rect 566 321 572 323
rect 566 319 568 321
rect 570 319 572 321
rect 566 317 572 319
rect 560 314 562 317
rect 570 314 572 317
rect 525 312 527 314
rect 529 312 531 314
rect 525 310 531 312
rect 529 307 531 310
rect 499 295 501 300
rect 509 295 511 300
rect 421 290 423 294
rect 428 290 430 294
rect 439 290 441 294
rect 461 290 463 294
rect 472 290 474 294
rect 479 290 481 294
rect 519 292 521 297
rect 550 303 552 308
rect 560 303 562 308
rect 598 312 600 325
rect 608 323 610 334
rect 670 351 672 356
rect 677 351 679 356
rect 695 354 697 358
rect 705 354 707 358
rect 715 354 717 358
rect 737 354 739 358
rect 747 354 749 358
rect 757 354 759 358
rect 660 342 662 347
rect 618 323 620 327
rect 604 321 610 323
rect 604 319 606 321
rect 608 319 610 321
rect 604 317 610 319
rect 614 321 620 323
rect 614 319 616 321
rect 618 319 620 321
rect 614 317 620 319
rect 605 312 607 317
rect 618 312 620 317
rect 647 316 649 329
rect 660 326 662 329
rect 775 351 777 356
rect 782 351 784 356
rect 805 354 807 358
rect 826 354 828 358
rect 833 354 835 358
rect 792 342 794 347
rect 924 354 926 358
rect 846 344 848 349
rect 874 347 876 352
rect 884 347 886 352
rect 826 330 828 333
rect 792 326 794 329
rect 653 324 662 326
rect 653 322 655 324
rect 657 322 659 324
rect 670 323 672 326
rect 677 323 679 326
rect 695 323 697 326
rect 705 323 707 326
rect 715 323 717 326
rect 737 323 739 326
rect 747 323 749 326
rect 757 323 759 326
rect 775 323 777 326
rect 782 323 784 326
rect 792 324 801 326
rect 653 320 659 322
rect 647 314 653 316
rect 647 312 649 314
rect 651 312 653 314
rect 570 300 572 305
rect 647 310 653 312
rect 647 307 649 310
rect 657 307 659 320
rect 667 321 673 323
rect 667 319 669 321
rect 671 319 673 321
rect 667 317 673 319
rect 677 321 699 323
rect 677 319 688 321
rect 690 319 695 321
rect 697 319 699 321
rect 677 317 699 319
rect 703 321 709 323
rect 703 319 705 321
rect 707 319 709 321
rect 703 317 709 319
rect 713 321 719 323
rect 713 319 715 321
rect 717 319 719 321
rect 713 317 719 319
rect 735 321 741 323
rect 735 319 737 321
rect 739 319 741 321
rect 735 317 741 319
rect 745 321 751 323
rect 745 319 747 321
rect 749 319 751 321
rect 745 317 751 319
rect 755 321 777 323
rect 755 319 757 321
rect 759 319 764 321
rect 766 319 777 321
rect 755 317 777 319
rect 781 321 787 323
rect 781 319 783 321
rect 785 319 787 321
rect 781 317 787 319
rect 667 314 669 317
rect 677 314 679 317
rect 697 314 699 317
rect 704 314 706 317
rect 598 296 600 301
rect 605 296 607 301
rect 529 290 531 294
rect 618 299 620 303
rect 647 290 649 294
rect 657 292 659 297
rect 667 295 669 300
rect 677 295 679 300
rect 715 308 717 317
rect 737 308 739 317
rect 748 314 750 317
rect 755 314 757 317
rect 775 314 777 317
rect 785 314 787 317
rect 795 322 797 324
rect 799 322 801 324
rect 795 320 801 322
rect 795 307 797 320
rect 805 316 807 329
rect 822 328 828 330
rect 822 326 824 328
rect 826 326 828 328
rect 822 324 828 326
rect 801 314 807 316
rect 826 314 828 324
rect 833 323 835 333
rect 894 345 896 349
rect 874 331 876 334
rect 870 329 876 331
rect 870 327 872 329
rect 874 327 876 329
rect 846 323 848 326
rect 870 325 876 327
rect 832 321 838 323
rect 832 319 834 321
rect 836 319 838 321
rect 832 317 838 319
rect 842 321 848 323
rect 842 319 844 321
rect 846 319 848 321
rect 842 317 848 319
rect 836 314 838 317
rect 846 314 848 317
rect 801 312 803 314
rect 805 312 807 314
rect 801 310 807 312
rect 805 307 807 310
rect 775 295 777 300
rect 785 295 787 300
rect 697 290 699 294
rect 704 290 706 294
rect 715 290 717 294
rect 737 290 739 294
rect 748 290 750 294
rect 755 290 757 294
rect 795 292 797 297
rect 826 303 828 308
rect 836 303 838 308
rect 874 312 876 325
rect 884 323 886 334
rect 947 351 949 356
rect 954 351 956 356
rect 972 354 974 358
rect 982 354 984 358
rect 992 354 994 358
rect 1014 354 1016 358
rect 1024 354 1026 358
rect 1034 354 1036 358
rect 937 342 939 347
rect 894 323 896 327
rect 880 321 886 323
rect 880 319 882 321
rect 884 319 886 321
rect 880 317 886 319
rect 890 321 896 323
rect 890 319 892 321
rect 894 319 896 321
rect 890 317 896 319
rect 881 312 883 317
rect 894 312 896 317
rect 924 316 926 329
rect 937 326 939 329
rect 1052 351 1054 356
rect 1059 351 1061 356
rect 1082 354 1084 358
rect 1103 354 1105 358
rect 1110 354 1112 358
rect 1069 342 1071 347
rect 1123 344 1125 349
rect 1103 330 1105 333
rect 1069 326 1071 329
rect 930 324 939 326
rect 930 322 932 324
rect 934 322 936 324
rect 947 323 949 326
rect 954 323 956 326
rect 972 323 974 326
rect 982 323 984 326
rect 992 323 994 326
rect 1014 323 1016 326
rect 1024 323 1026 326
rect 1034 323 1036 326
rect 1052 323 1054 326
rect 1059 323 1061 326
rect 1069 324 1078 326
rect 930 320 936 322
rect 924 314 930 316
rect 924 312 926 314
rect 928 312 930 314
rect 846 300 848 305
rect 924 310 930 312
rect 924 307 926 310
rect 934 307 936 320
rect 944 321 950 323
rect 944 319 946 321
rect 948 319 950 321
rect 944 317 950 319
rect 954 321 976 323
rect 954 319 965 321
rect 967 319 972 321
rect 974 319 976 321
rect 954 317 976 319
rect 980 321 986 323
rect 980 319 982 321
rect 984 319 986 321
rect 980 317 986 319
rect 990 321 996 323
rect 990 319 992 321
rect 994 319 996 321
rect 990 317 996 319
rect 1012 321 1018 323
rect 1012 319 1014 321
rect 1016 319 1018 321
rect 1012 317 1018 319
rect 1022 321 1028 323
rect 1022 319 1024 321
rect 1026 319 1028 321
rect 1022 317 1028 319
rect 1032 321 1054 323
rect 1032 319 1034 321
rect 1036 319 1041 321
rect 1043 319 1054 321
rect 1032 317 1054 319
rect 1058 321 1064 323
rect 1058 319 1060 321
rect 1062 319 1064 321
rect 1058 317 1064 319
rect 944 314 946 317
rect 954 314 956 317
rect 974 314 976 317
rect 981 314 983 317
rect 874 296 876 301
rect 881 296 883 301
rect 805 290 807 294
rect 894 299 896 303
rect 924 290 926 294
rect 934 292 936 297
rect 944 295 946 300
rect 954 295 956 300
rect 992 308 994 317
rect 1014 308 1016 317
rect 1025 314 1027 317
rect 1032 314 1034 317
rect 1052 314 1054 317
rect 1062 314 1064 317
rect 1072 322 1074 324
rect 1076 322 1078 324
rect 1072 320 1078 322
rect 1072 307 1074 320
rect 1082 316 1084 329
rect 1099 328 1105 330
rect 1099 326 1101 328
rect 1103 326 1105 328
rect 1099 324 1105 326
rect 1078 314 1084 316
rect 1103 314 1105 324
rect 1110 323 1112 333
rect 1123 323 1125 326
rect 1109 321 1115 323
rect 1109 319 1111 321
rect 1113 319 1115 321
rect 1109 317 1115 319
rect 1119 321 1125 323
rect 1119 319 1121 321
rect 1123 319 1125 321
rect 1119 317 1125 319
rect 1113 314 1115 317
rect 1123 314 1125 317
rect 1078 312 1080 314
rect 1082 312 1084 314
rect 1078 310 1084 312
rect 1082 307 1084 310
rect 1052 295 1054 300
rect 1062 295 1064 300
rect 974 290 976 294
rect 981 290 983 294
rect 992 290 994 294
rect 1014 290 1016 294
rect 1025 290 1027 294
rect 1032 290 1034 294
rect 1072 292 1074 297
rect 1103 303 1105 308
rect 1113 303 1115 308
rect 1123 300 1125 305
rect 1082 290 1084 294
rect -273 284 -248 286
rect -273 276 -271 284
rect -260 276 -258 280
rect -250 276 -248 284
rect -240 279 -238 284
rect -233 279 -231 284
rect -208 282 -206 286
rect -276 274 -271 276
rect -276 271 -274 274
rect -198 279 -196 284
rect -158 282 -156 286
rect -151 282 -149 286
rect -140 282 -138 286
rect -118 282 -116 286
rect -107 282 -105 286
rect -100 282 -98 286
rect -188 276 -186 281
rect -178 276 -176 281
rect -260 264 -258 267
rect -267 262 -258 264
rect -250 263 -248 267
rect -240 264 -238 267
rect -276 254 -274 262
rect -267 260 -265 262
rect -263 260 -258 262
rect -267 258 -258 260
rect -242 262 -238 264
rect -242 259 -240 262
rect -260 254 -258 258
rect -246 257 -240 259
rect -233 258 -231 267
rect -208 266 -206 269
rect -208 264 -202 266
rect -208 262 -206 264
rect -204 262 -202 264
rect -208 260 -202 262
rect -246 255 -244 257
rect -242 255 -240 257
rect -279 252 -266 254
rect -260 252 -250 254
rect -246 253 -240 255
rect -279 251 -277 252
rect -283 249 -277 251
rect -268 249 -266 252
rect -252 249 -250 252
rect -242 249 -240 253
rect -236 256 -230 258
rect -236 254 -234 256
rect -232 254 -230 256
rect -236 252 -230 254
rect -232 249 -230 252
rect -283 247 -281 249
rect -279 247 -277 249
rect -283 245 -277 247
rect -252 227 -250 231
rect -242 227 -240 231
rect -268 218 -266 222
rect -208 247 -206 260
rect -198 256 -196 269
rect -202 254 -196 256
rect -202 252 -200 254
rect -198 252 -196 254
rect -188 259 -186 262
rect -178 259 -176 262
rect -158 259 -156 262
rect -151 259 -149 262
rect -140 259 -138 268
rect -118 259 -116 268
rect -80 276 -78 281
rect -70 276 -68 281
rect -60 279 -58 284
rect -50 282 -48 286
rect -107 259 -105 262
rect -100 259 -98 262
rect -80 259 -78 262
rect -70 259 -68 262
rect -188 257 -182 259
rect -188 255 -186 257
rect -184 255 -182 257
rect -188 253 -182 255
rect -178 257 -156 259
rect -178 255 -167 257
rect -165 255 -160 257
rect -158 255 -156 257
rect -178 253 -156 255
rect -152 257 -146 259
rect -152 255 -150 257
rect -148 255 -146 257
rect -152 253 -146 255
rect -142 257 -136 259
rect -142 255 -140 257
rect -138 255 -136 257
rect -142 253 -136 255
rect -120 257 -114 259
rect -120 255 -118 257
rect -116 255 -114 257
rect -120 253 -114 255
rect -110 257 -104 259
rect -110 255 -108 257
rect -106 255 -104 257
rect -110 253 -104 255
rect -100 257 -78 259
rect -100 255 -98 257
rect -96 255 -91 257
rect -89 255 -78 257
rect -100 253 -78 255
rect -74 257 -68 259
rect -74 255 -72 257
rect -70 255 -68 257
rect -74 253 -68 255
rect -60 256 -58 269
rect -50 266 -48 269
rect -54 264 -48 266
rect -54 262 -52 264
rect -50 262 -48 264
rect -29 268 -27 273
rect -19 268 -17 273
rect -9 271 -7 276
rect 14 275 16 280
rect 21 275 23 280
rect 34 273 36 277
rect 54 275 56 280
rect 61 275 63 280
rect 94 282 96 286
rect 74 273 76 277
rect 104 279 106 284
rect 144 282 146 286
rect 151 282 153 286
rect 162 282 164 286
rect 184 282 186 286
rect 195 282 197 286
rect 202 282 204 286
rect 114 276 116 281
rect 124 276 126 281
rect 94 266 96 269
rect 94 264 100 266
rect -54 260 -48 262
rect -60 254 -54 256
rect -202 250 -193 252
rect -185 250 -183 253
rect -178 250 -176 253
rect -160 250 -158 253
rect -150 250 -148 253
rect -140 250 -138 253
rect -118 250 -116 253
rect -108 250 -106 253
rect -98 250 -96 253
rect -80 250 -78 253
rect -73 250 -71 253
rect -60 252 -58 254
rect -56 252 -54 254
rect -63 250 -54 252
rect -195 247 -193 250
rect -195 229 -193 234
rect -232 218 -230 222
rect -208 218 -206 222
rect -185 220 -183 225
rect -178 220 -176 225
rect -63 247 -61 250
rect -50 247 -48 260
rect -29 252 -27 262
rect -19 259 -17 262
rect -9 259 -7 262
rect -23 257 -17 259
rect -23 255 -21 257
rect -19 255 -17 257
rect -23 253 -17 255
rect -13 257 -7 259
rect -13 255 -11 257
rect -9 255 -7 257
rect -13 253 -7 255
rect -33 250 -27 252
rect -33 248 -31 250
rect -29 248 -27 250
rect -63 229 -61 234
rect -160 218 -158 222
rect -150 218 -148 222
rect -140 218 -138 222
rect -118 218 -116 222
rect -108 218 -106 222
rect -98 218 -96 222
rect -80 220 -78 225
rect -73 220 -71 225
rect -33 246 -27 248
rect -29 243 -27 246
rect -22 243 -20 253
rect -9 250 -7 253
rect 14 251 16 264
rect 21 259 23 264
rect 34 259 36 264
rect 20 257 26 259
rect 20 255 22 257
rect 24 255 26 257
rect 20 253 26 255
rect 30 257 36 259
rect 30 255 32 257
rect 34 255 36 257
rect 30 253 36 255
rect 10 249 16 251
rect 10 247 12 249
rect 14 247 16 249
rect 10 245 16 247
rect 14 242 16 245
rect 24 242 26 253
rect 34 249 36 253
rect 54 251 56 264
rect 61 259 63 264
rect 74 259 76 264
rect 60 257 66 259
rect 60 255 62 257
rect 64 255 66 257
rect 60 253 66 255
rect 70 257 76 259
rect 70 255 72 257
rect 74 255 76 257
rect 70 253 76 255
rect 50 249 56 251
rect -9 227 -7 232
rect 50 247 52 249
rect 54 247 56 249
rect 50 245 56 247
rect 54 242 56 245
rect 64 242 66 253
rect 74 249 76 253
rect 94 262 96 264
rect 98 262 100 264
rect 94 260 100 262
rect 14 224 16 229
rect 24 224 26 229
rect 34 227 36 231
rect 94 247 96 260
rect 104 256 106 269
rect 100 254 106 256
rect 100 252 102 254
rect 104 252 106 254
rect 114 259 116 262
rect 124 259 126 262
rect 144 259 146 262
rect 151 259 153 262
rect 162 259 164 268
rect 184 259 186 268
rect 222 276 224 281
rect 232 276 234 281
rect 242 279 244 284
rect 252 282 254 286
rect 195 259 197 262
rect 202 259 204 262
rect 222 259 224 262
rect 232 259 234 262
rect 114 257 120 259
rect 114 255 116 257
rect 118 255 120 257
rect 114 253 120 255
rect 124 257 146 259
rect 124 255 135 257
rect 137 255 142 257
rect 144 255 146 257
rect 124 253 146 255
rect 150 257 156 259
rect 150 255 152 257
rect 154 255 156 257
rect 150 253 156 255
rect 160 257 166 259
rect 160 255 162 257
rect 164 255 166 257
rect 160 253 166 255
rect 182 257 188 259
rect 182 255 184 257
rect 186 255 188 257
rect 182 253 188 255
rect 192 257 198 259
rect 192 255 194 257
rect 196 255 198 257
rect 192 253 198 255
rect 202 257 224 259
rect 202 255 204 257
rect 206 255 211 257
rect 213 255 224 257
rect 202 253 224 255
rect 228 257 234 259
rect 228 255 230 257
rect 232 255 234 257
rect 228 253 234 255
rect 242 256 244 269
rect 252 266 254 269
rect 248 264 254 266
rect 248 262 250 264
rect 252 262 254 264
rect 273 268 275 273
rect 283 268 285 273
rect 293 271 295 276
rect 321 275 323 280
rect 328 275 330 280
rect 371 282 373 286
rect 341 273 343 277
rect 381 279 383 284
rect 421 282 423 286
rect 428 282 430 286
rect 439 282 441 286
rect 461 282 463 286
rect 472 282 474 286
rect 479 282 481 286
rect 391 276 393 281
rect 401 276 403 281
rect 371 266 373 269
rect 371 264 377 266
rect 248 260 254 262
rect 242 254 248 256
rect 100 250 109 252
rect 117 250 119 253
rect 124 250 126 253
rect 142 250 144 253
rect 152 250 154 253
rect 162 250 164 253
rect 184 250 186 253
rect 194 250 196 253
rect 204 250 206 253
rect 222 250 224 253
rect 229 250 231 253
rect 242 252 244 254
rect 246 252 248 254
rect 239 250 248 252
rect 107 247 109 250
rect -50 218 -48 222
rect -29 218 -27 222
rect -22 218 -20 222
rect 54 224 56 229
rect 64 224 66 229
rect 74 227 76 231
rect 107 229 109 234
rect 94 218 96 222
rect 117 220 119 225
rect 124 220 126 225
rect 239 247 241 250
rect 252 247 254 260
rect 273 252 275 262
rect 283 259 285 262
rect 293 259 295 262
rect 279 257 285 259
rect 279 255 281 257
rect 283 255 285 257
rect 279 253 285 255
rect 289 257 295 259
rect 289 255 291 257
rect 293 255 295 257
rect 289 253 295 255
rect 269 250 275 252
rect 269 248 271 250
rect 273 248 275 250
rect 239 229 241 234
rect 142 218 144 222
rect 152 218 154 222
rect 162 218 164 222
rect 184 218 186 222
rect 194 218 196 222
rect 204 218 206 222
rect 222 220 224 225
rect 229 220 231 225
rect 269 246 275 248
rect 273 243 275 246
rect 280 243 282 253
rect 293 250 295 253
rect 321 251 323 264
rect 328 259 330 264
rect 341 259 343 264
rect 327 257 333 259
rect 327 255 329 257
rect 331 255 333 257
rect 327 253 333 255
rect 337 257 343 259
rect 337 255 339 257
rect 341 255 343 257
rect 337 253 343 255
rect 317 249 323 251
rect 317 247 319 249
rect 321 247 323 249
rect 317 245 323 247
rect 321 242 323 245
rect 331 242 333 253
rect 341 249 343 253
rect 371 262 373 264
rect 375 262 377 264
rect 371 260 377 262
rect 293 227 295 232
rect 371 247 373 260
rect 381 256 383 269
rect 377 254 383 256
rect 377 252 379 254
rect 381 252 383 254
rect 391 259 393 262
rect 401 259 403 262
rect 421 259 423 262
rect 428 259 430 262
rect 439 259 441 268
rect 461 259 463 268
rect 499 276 501 281
rect 509 276 511 281
rect 519 279 521 284
rect 529 282 531 286
rect 472 259 474 262
rect 479 259 481 262
rect 499 259 501 262
rect 509 259 511 262
rect 391 257 397 259
rect 391 255 393 257
rect 395 255 397 257
rect 391 253 397 255
rect 401 257 423 259
rect 401 255 412 257
rect 414 255 419 257
rect 421 255 423 257
rect 401 253 423 255
rect 427 257 433 259
rect 427 255 429 257
rect 431 255 433 257
rect 427 253 433 255
rect 437 257 443 259
rect 437 255 439 257
rect 441 255 443 257
rect 437 253 443 255
rect 459 257 465 259
rect 459 255 461 257
rect 463 255 465 257
rect 459 253 465 255
rect 469 257 475 259
rect 469 255 471 257
rect 473 255 475 257
rect 469 253 475 255
rect 479 257 501 259
rect 479 255 481 257
rect 483 255 488 257
rect 490 255 501 257
rect 479 253 501 255
rect 505 257 511 259
rect 505 255 507 257
rect 509 255 511 257
rect 505 253 511 255
rect 519 256 521 269
rect 529 266 531 269
rect 525 264 531 266
rect 525 262 527 264
rect 529 262 531 264
rect 550 268 552 273
rect 560 268 562 273
rect 570 271 572 276
rect 598 275 600 280
rect 605 275 607 280
rect 647 282 649 286
rect 618 273 620 277
rect 657 279 659 284
rect 697 282 699 286
rect 704 282 706 286
rect 715 282 717 286
rect 737 282 739 286
rect 748 282 750 286
rect 755 282 757 286
rect 667 276 669 281
rect 677 276 679 281
rect 647 266 649 269
rect 647 264 653 266
rect 525 260 531 262
rect 519 254 525 256
rect 377 250 386 252
rect 394 250 396 253
rect 401 250 403 253
rect 419 250 421 253
rect 429 250 431 253
rect 439 250 441 253
rect 461 250 463 253
rect 471 250 473 253
rect 481 250 483 253
rect 499 250 501 253
rect 506 250 508 253
rect 519 252 521 254
rect 523 252 525 254
rect 516 250 525 252
rect 384 247 386 250
rect 321 224 323 229
rect 331 224 333 229
rect 341 227 343 231
rect 252 218 254 222
rect 273 218 275 222
rect 280 218 282 222
rect 384 229 386 234
rect 371 218 373 222
rect 394 220 396 225
rect 401 220 403 225
rect 516 247 518 250
rect 529 247 531 260
rect 550 252 552 262
rect 560 259 562 262
rect 570 259 572 262
rect 556 257 562 259
rect 556 255 558 257
rect 560 255 562 257
rect 556 253 562 255
rect 566 257 572 259
rect 566 255 568 257
rect 570 255 572 257
rect 566 253 572 255
rect 546 250 552 252
rect 546 248 548 250
rect 550 248 552 250
rect 516 229 518 234
rect 419 218 421 222
rect 429 218 431 222
rect 439 218 441 222
rect 461 218 463 222
rect 471 218 473 222
rect 481 218 483 222
rect 499 220 501 225
rect 506 220 508 225
rect 546 246 552 248
rect 550 243 552 246
rect 557 243 559 253
rect 570 250 572 253
rect 598 251 600 264
rect 605 259 607 264
rect 618 259 620 264
rect 604 257 610 259
rect 604 255 606 257
rect 608 255 610 257
rect 604 253 610 255
rect 614 257 620 259
rect 614 255 616 257
rect 618 255 620 257
rect 614 253 620 255
rect 594 249 600 251
rect 594 247 596 249
rect 598 247 600 249
rect 594 245 600 247
rect 598 242 600 245
rect 608 242 610 253
rect 618 249 620 253
rect 647 262 649 264
rect 651 262 653 264
rect 647 260 653 262
rect 570 227 572 232
rect 647 247 649 260
rect 657 256 659 269
rect 653 254 659 256
rect 653 252 655 254
rect 657 252 659 254
rect 667 259 669 262
rect 677 259 679 262
rect 697 259 699 262
rect 704 259 706 262
rect 715 259 717 268
rect 737 259 739 268
rect 775 276 777 281
rect 785 276 787 281
rect 795 279 797 284
rect 805 282 807 286
rect 748 259 750 262
rect 755 259 757 262
rect 775 259 777 262
rect 785 259 787 262
rect 667 257 673 259
rect 667 255 669 257
rect 671 255 673 257
rect 667 253 673 255
rect 677 257 699 259
rect 677 255 688 257
rect 690 255 695 257
rect 697 255 699 257
rect 677 253 699 255
rect 703 257 709 259
rect 703 255 705 257
rect 707 255 709 257
rect 703 253 709 255
rect 713 257 719 259
rect 713 255 715 257
rect 717 255 719 257
rect 713 253 719 255
rect 735 257 741 259
rect 735 255 737 257
rect 739 255 741 257
rect 735 253 741 255
rect 745 257 751 259
rect 745 255 747 257
rect 749 255 751 257
rect 745 253 751 255
rect 755 257 777 259
rect 755 255 757 257
rect 759 255 764 257
rect 766 255 777 257
rect 755 253 777 255
rect 781 257 787 259
rect 781 255 783 257
rect 785 255 787 257
rect 781 253 787 255
rect 795 256 797 269
rect 805 266 807 269
rect 801 264 807 266
rect 801 262 803 264
rect 805 262 807 264
rect 826 268 828 273
rect 836 268 838 273
rect 846 271 848 276
rect 874 275 876 280
rect 881 275 883 280
rect 924 282 926 286
rect 894 273 896 277
rect 934 279 936 284
rect 974 282 976 286
rect 981 282 983 286
rect 992 282 994 286
rect 1014 282 1016 286
rect 1025 282 1027 286
rect 1032 282 1034 286
rect 944 276 946 281
rect 954 276 956 281
rect 924 266 926 269
rect 924 264 930 266
rect 801 260 807 262
rect 795 254 801 256
rect 653 250 662 252
rect 670 250 672 253
rect 677 250 679 253
rect 695 250 697 253
rect 705 250 707 253
rect 715 250 717 253
rect 737 250 739 253
rect 747 250 749 253
rect 757 250 759 253
rect 775 250 777 253
rect 782 250 784 253
rect 795 252 797 254
rect 799 252 801 254
rect 792 250 801 252
rect 660 247 662 250
rect 598 224 600 229
rect 608 224 610 229
rect 618 227 620 231
rect 529 218 531 222
rect 550 218 552 222
rect 557 218 559 222
rect 660 229 662 234
rect 647 218 649 222
rect 670 220 672 225
rect 677 220 679 225
rect 792 247 794 250
rect 805 247 807 260
rect 826 252 828 262
rect 836 259 838 262
rect 846 259 848 262
rect 832 257 838 259
rect 832 255 834 257
rect 836 255 838 257
rect 832 253 838 255
rect 842 257 848 259
rect 842 255 844 257
rect 846 255 848 257
rect 842 253 848 255
rect 822 250 828 252
rect 822 248 824 250
rect 826 248 828 250
rect 792 229 794 234
rect 695 218 697 222
rect 705 218 707 222
rect 715 218 717 222
rect 737 218 739 222
rect 747 218 749 222
rect 757 218 759 222
rect 775 220 777 225
rect 782 220 784 225
rect 822 246 828 248
rect 826 243 828 246
rect 833 243 835 253
rect 846 250 848 253
rect 874 251 876 264
rect 881 259 883 264
rect 894 259 896 264
rect 880 257 886 259
rect 880 255 882 257
rect 884 255 886 257
rect 880 253 886 255
rect 890 257 896 259
rect 890 255 892 257
rect 894 255 896 257
rect 890 253 896 255
rect 870 249 876 251
rect 870 247 872 249
rect 874 247 876 249
rect 870 245 876 247
rect 874 242 876 245
rect 884 242 886 253
rect 894 249 896 253
rect 924 262 926 264
rect 928 262 930 264
rect 924 260 930 262
rect 846 227 848 232
rect 924 247 926 260
rect 934 256 936 269
rect 930 254 936 256
rect 930 252 932 254
rect 934 252 936 254
rect 944 259 946 262
rect 954 259 956 262
rect 974 259 976 262
rect 981 259 983 262
rect 992 259 994 268
rect 1014 259 1016 268
rect 1052 276 1054 281
rect 1062 276 1064 281
rect 1072 279 1074 284
rect 1082 282 1084 286
rect 1025 259 1027 262
rect 1032 259 1034 262
rect 1052 259 1054 262
rect 1062 259 1064 262
rect 944 257 950 259
rect 944 255 946 257
rect 948 255 950 257
rect 944 253 950 255
rect 954 257 976 259
rect 954 255 965 257
rect 967 255 972 257
rect 974 255 976 257
rect 954 253 976 255
rect 980 257 986 259
rect 980 255 982 257
rect 984 255 986 257
rect 980 253 986 255
rect 990 257 996 259
rect 990 255 992 257
rect 994 255 996 257
rect 990 253 996 255
rect 1012 257 1018 259
rect 1012 255 1014 257
rect 1016 255 1018 257
rect 1012 253 1018 255
rect 1022 257 1028 259
rect 1022 255 1024 257
rect 1026 255 1028 257
rect 1022 253 1028 255
rect 1032 257 1054 259
rect 1032 255 1034 257
rect 1036 255 1041 257
rect 1043 255 1054 257
rect 1032 253 1054 255
rect 1058 257 1064 259
rect 1058 255 1060 257
rect 1062 255 1064 257
rect 1058 253 1064 255
rect 1072 256 1074 269
rect 1082 266 1084 269
rect 1078 264 1084 266
rect 1078 262 1080 264
rect 1082 262 1084 264
rect 1103 268 1105 273
rect 1113 268 1115 273
rect 1123 271 1125 276
rect 1078 260 1084 262
rect 1072 254 1078 256
rect 930 250 939 252
rect 947 250 949 253
rect 954 250 956 253
rect 972 250 974 253
rect 982 250 984 253
rect 992 250 994 253
rect 1014 250 1016 253
rect 1024 250 1026 253
rect 1034 250 1036 253
rect 1052 250 1054 253
rect 1059 250 1061 253
rect 1072 252 1074 254
rect 1076 252 1078 254
rect 1069 250 1078 252
rect 937 247 939 250
rect 874 224 876 229
rect 884 224 886 229
rect 894 227 896 231
rect 805 218 807 222
rect 826 218 828 222
rect 833 218 835 222
rect 937 229 939 234
rect 924 218 926 222
rect 947 220 949 225
rect 954 220 956 225
rect 1069 247 1071 250
rect 1082 247 1084 260
rect 1103 252 1105 262
rect 1113 259 1115 262
rect 1123 259 1125 262
rect 1109 257 1115 259
rect 1109 255 1111 257
rect 1113 255 1115 257
rect 1109 253 1115 255
rect 1119 257 1125 259
rect 1119 255 1121 257
rect 1123 255 1125 257
rect 1119 253 1125 255
rect 1099 250 1105 252
rect 1099 248 1101 250
rect 1103 248 1105 250
rect 1069 229 1071 234
rect 972 218 974 222
rect 982 218 984 222
rect 992 218 994 222
rect 1014 218 1016 222
rect 1024 218 1026 222
rect 1034 218 1036 222
rect 1052 220 1054 225
rect 1059 220 1061 225
rect 1099 246 1105 248
rect 1103 243 1105 246
rect 1110 243 1112 253
rect 1123 250 1125 253
rect 1123 227 1125 232
rect 1082 218 1084 222
rect 1103 218 1105 222
rect 1110 218 1112 222
rect -268 210 -266 214
rect -283 185 -277 187
rect -283 183 -281 185
rect -279 183 -277 185
rect -232 210 -230 214
rect -208 210 -206 214
rect -252 201 -250 205
rect -242 201 -240 205
rect -185 207 -183 212
rect -178 207 -176 212
rect -160 210 -158 214
rect -150 210 -148 214
rect -140 210 -138 214
rect -118 210 -116 214
rect -108 210 -106 214
rect -98 210 -96 214
rect -195 198 -193 203
rect -283 181 -277 183
rect -279 180 -277 181
rect -268 180 -266 183
rect -252 180 -250 183
rect -279 178 -266 180
rect -260 178 -250 180
rect -242 179 -240 183
rect -232 180 -230 183
rect -276 170 -274 178
rect -260 174 -258 178
rect -267 172 -258 174
rect -246 177 -240 179
rect -246 175 -244 177
rect -242 175 -240 177
rect -246 173 -240 175
rect -236 178 -230 180
rect -236 176 -234 178
rect -232 176 -230 178
rect -236 174 -230 176
rect -267 170 -265 172
rect -263 170 -258 172
rect -267 168 -258 170
rect -242 170 -240 173
rect -260 165 -258 168
rect -250 165 -248 169
rect -242 168 -238 170
rect -240 165 -238 168
rect -233 165 -231 174
rect -208 172 -206 185
rect -195 182 -193 185
rect -80 207 -78 212
rect -73 207 -71 212
rect -50 210 -48 214
rect -29 210 -27 214
rect -22 210 -20 214
rect -63 198 -61 203
rect -9 200 -7 205
rect 14 203 16 208
rect 24 203 26 208
rect 94 210 96 214
rect -29 186 -27 189
rect -63 182 -61 185
rect -202 180 -193 182
rect -202 178 -200 180
rect -198 178 -196 180
rect -185 179 -183 182
rect -178 179 -176 182
rect -160 179 -158 182
rect -150 179 -148 182
rect -140 179 -138 182
rect -118 179 -116 182
rect -108 179 -106 182
rect -98 179 -96 182
rect -80 179 -78 182
rect -73 179 -71 182
rect -63 180 -54 182
rect -202 176 -196 178
rect -208 170 -202 172
rect -208 168 -206 170
rect -204 168 -202 170
rect -208 166 -202 168
rect -276 158 -274 161
rect -276 156 -271 158
rect -273 148 -271 156
rect -260 152 -258 156
rect -250 148 -248 156
rect -208 163 -206 166
rect -198 163 -196 176
rect -188 177 -182 179
rect -188 175 -186 177
rect -184 175 -182 177
rect -188 173 -182 175
rect -178 177 -156 179
rect -178 175 -167 177
rect -165 175 -160 177
rect -158 175 -156 177
rect -178 173 -156 175
rect -152 177 -146 179
rect -152 175 -150 177
rect -148 175 -146 177
rect -152 173 -146 175
rect -142 177 -136 179
rect -142 175 -140 177
rect -138 175 -136 177
rect -142 173 -136 175
rect -120 177 -114 179
rect -120 175 -118 177
rect -116 175 -114 177
rect -120 173 -114 175
rect -110 177 -104 179
rect -110 175 -108 177
rect -106 175 -104 177
rect -110 173 -104 175
rect -100 177 -78 179
rect -100 175 -98 177
rect -96 175 -91 177
rect -89 175 -78 177
rect -100 173 -78 175
rect -74 177 -68 179
rect -74 175 -72 177
rect -70 175 -68 177
rect -74 173 -68 175
rect -188 170 -186 173
rect -178 170 -176 173
rect -158 170 -156 173
rect -151 170 -149 173
rect -240 148 -238 153
rect -233 148 -231 153
rect -273 146 -248 148
rect -208 146 -206 150
rect -198 148 -196 153
rect -188 151 -186 156
rect -178 151 -176 156
rect -140 164 -138 173
rect -118 164 -116 173
rect -107 170 -105 173
rect -100 170 -98 173
rect -80 170 -78 173
rect -70 170 -68 173
rect -60 178 -58 180
rect -56 178 -54 180
rect -60 176 -54 178
rect -60 163 -58 176
rect -50 172 -48 185
rect -33 184 -27 186
rect -33 182 -31 184
rect -29 182 -27 184
rect -33 180 -27 182
rect -54 170 -48 172
rect -29 170 -27 180
rect -22 179 -20 189
rect 34 201 36 205
rect 54 203 56 208
rect 64 203 66 208
rect 14 187 16 190
rect 10 185 16 187
rect 10 183 12 185
rect 14 183 16 185
rect -9 179 -7 182
rect 10 181 16 183
rect -23 177 -17 179
rect -23 175 -21 177
rect -19 175 -17 177
rect -23 173 -17 175
rect -13 177 -7 179
rect -13 175 -11 177
rect -9 175 -7 177
rect -13 173 -7 175
rect -19 170 -17 173
rect -9 170 -7 173
rect -54 168 -52 170
rect -50 168 -48 170
rect -54 166 -48 168
rect -50 163 -48 166
rect -80 151 -78 156
rect -70 151 -68 156
rect -158 146 -156 150
rect -151 146 -149 150
rect -140 146 -138 150
rect -118 146 -116 150
rect -107 146 -105 150
rect -100 146 -98 150
rect -60 148 -58 153
rect -29 159 -27 164
rect -19 159 -17 164
rect 14 168 16 181
rect 24 179 26 190
rect 74 201 76 205
rect 54 187 56 190
rect 50 185 56 187
rect 50 183 52 185
rect 54 183 56 185
rect 34 179 36 183
rect 50 181 56 183
rect 20 177 26 179
rect 20 175 22 177
rect 24 175 26 177
rect 20 173 26 175
rect 30 177 36 179
rect 30 175 32 177
rect 34 175 36 177
rect 30 173 36 175
rect 21 168 23 173
rect 34 168 36 173
rect 54 168 56 181
rect 64 179 66 190
rect 117 207 119 212
rect 124 207 126 212
rect 142 210 144 214
rect 152 210 154 214
rect 162 210 164 214
rect 184 210 186 214
rect 194 210 196 214
rect 204 210 206 214
rect 107 198 109 203
rect 74 179 76 183
rect 60 177 66 179
rect 60 175 62 177
rect 64 175 66 177
rect 60 173 66 175
rect 70 177 76 179
rect 70 175 72 177
rect 74 175 76 177
rect 70 173 76 175
rect 61 168 63 173
rect 74 168 76 173
rect 94 172 96 185
rect 107 182 109 185
rect 222 207 224 212
rect 229 207 231 212
rect 252 210 254 214
rect 273 210 275 214
rect 280 210 282 214
rect 239 198 241 203
rect 371 210 373 214
rect 293 200 295 205
rect 321 203 323 208
rect 331 203 333 208
rect 273 186 275 189
rect 239 182 241 185
rect 100 180 109 182
rect 100 178 102 180
rect 104 178 106 180
rect 117 179 119 182
rect 124 179 126 182
rect 142 179 144 182
rect 152 179 154 182
rect 162 179 164 182
rect 184 179 186 182
rect 194 179 196 182
rect 204 179 206 182
rect 222 179 224 182
rect 229 179 231 182
rect 239 180 248 182
rect 100 176 106 178
rect 94 170 100 172
rect 94 168 96 170
rect 98 168 100 170
rect -9 156 -7 161
rect 14 152 16 157
rect 21 152 23 157
rect -50 146 -48 150
rect 34 155 36 159
rect 94 166 100 168
rect 94 163 96 166
rect 104 163 106 176
rect 114 177 120 179
rect 114 175 116 177
rect 118 175 120 177
rect 114 173 120 175
rect 124 177 146 179
rect 124 175 135 177
rect 137 175 142 177
rect 144 175 146 177
rect 124 173 146 175
rect 150 177 156 179
rect 150 175 152 177
rect 154 175 156 177
rect 150 173 156 175
rect 160 177 166 179
rect 160 175 162 177
rect 164 175 166 177
rect 160 173 166 175
rect 182 177 188 179
rect 182 175 184 177
rect 186 175 188 177
rect 182 173 188 175
rect 192 177 198 179
rect 192 175 194 177
rect 196 175 198 177
rect 192 173 198 175
rect 202 177 224 179
rect 202 175 204 177
rect 206 175 211 177
rect 213 175 224 177
rect 202 173 224 175
rect 228 177 234 179
rect 228 175 230 177
rect 232 175 234 177
rect 228 173 234 175
rect 114 170 116 173
rect 124 170 126 173
rect 144 170 146 173
rect 151 170 153 173
rect 54 152 56 157
rect 61 152 63 157
rect 74 155 76 159
rect 94 146 96 150
rect 104 148 106 153
rect 114 151 116 156
rect 124 151 126 156
rect 162 164 164 173
rect 184 164 186 173
rect 195 170 197 173
rect 202 170 204 173
rect 222 170 224 173
rect 232 170 234 173
rect 242 178 244 180
rect 246 178 248 180
rect 242 176 248 178
rect 242 163 244 176
rect 252 172 254 185
rect 269 184 275 186
rect 269 182 271 184
rect 273 182 275 184
rect 269 180 275 182
rect 248 170 254 172
rect 273 170 275 180
rect 280 179 282 189
rect 341 201 343 205
rect 321 187 323 190
rect 317 185 323 187
rect 317 183 319 185
rect 321 183 323 185
rect 293 179 295 182
rect 317 181 323 183
rect 279 177 285 179
rect 279 175 281 177
rect 283 175 285 177
rect 279 173 285 175
rect 289 177 295 179
rect 289 175 291 177
rect 293 175 295 177
rect 289 173 295 175
rect 283 170 285 173
rect 293 170 295 173
rect 248 168 250 170
rect 252 168 254 170
rect 248 166 254 168
rect 252 163 254 166
rect 222 151 224 156
rect 232 151 234 156
rect 144 146 146 150
rect 151 146 153 150
rect 162 146 164 150
rect 184 146 186 150
rect 195 146 197 150
rect 202 146 204 150
rect 242 148 244 153
rect 273 159 275 164
rect 283 159 285 164
rect 321 168 323 181
rect 331 179 333 190
rect 394 207 396 212
rect 401 207 403 212
rect 419 210 421 214
rect 429 210 431 214
rect 439 210 441 214
rect 461 210 463 214
rect 471 210 473 214
rect 481 210 483 214
rect 384 198 386 203
rect 341 179 343 183
rect 327 177 333 179
rect 327 175 329 177
rect 331 175 333 177
rect 327 173 333 175
rect 337 177 343 179
rect 337 175 339 177
rect 341 175 343 177
rect 337 173 343 175
rect 328 168 330 173
rect 341 168 343 173
rect 371 172 373 185
rect 384 182 386 185
rect 499 207 501 212
rect 506 207 508 212
rect 529 210 531 214
rect 550 210 552 214
rect 557 210 559 214
rect 516 198 518 203
rect 647 210 649 214
rect 570 200 572 205
rect 598 203 600 208
rect 608 203 610 208
rect 550 186 552 189
rect 516 182 518 185
rect 377 180 386 182
rect 377 178 379 180
rect 381 178 383 180
rect 394 179 396 182
rect 401 179 403 182
rect 419 179 421 182
rect 429 179 431 182
rect 439 179 441 182
rect 461 179 463 182
rect 471 179 473 182
rect 481 179 483 182
rect 499 179 501 182
rect 506 179 508 182
rect 516 180 525 182
rect 377 176 383 178
rect 371 170 377 172
rect 371 168 373 170
rect 375 168 377 170
rect 293 156 295 161
rect 371 166 377 168
rect 371 163 373 166
rect 381 163 383 176
rect 391 177 397 179
rect 391 175 393 177
rect 395 175 397 177
rect 391 173 397 175
rect 401 177 423 179
rect 401 175 412 177
rect 414 175 419 177
rect 421 175 423 177
rect 401 173 423 175
rect 427 177 433 179
rect 427 175 429 177
rect 431 175 433 177
rect 427 173 433 175
rect 437 177 443 179
rect 437 175 439 177
rect 441 175 443 177
rect 437 173 443 175
rect 459 177 465 179
rect 459 175 461 177
rect 463 175 465 177
rect 459 173 465 175
rect 469 177 475 179
rect 469 175 471 177
rect 473 175 475 177
rect 469 173 475 175
rect 479 177 501 179
rect 479 175 481 177
rect 483 175 488 177
rect 490 175 501 177
rect 479 173 501 175
rect 505 177 511 179
rect 505 175 507 177
rect 509 175 511 177
rect 505 173 511 175
rect 391 170 393 173
rect 401 170 403 173
rect 421 170 423 173
rect 428 170 430 173
rect 321 152 323 157
rect 328 152 330 157
rect 252 146 254 150
rect 341 155 343 159
rect 371 146 373 150
rect 381 148 383 153
rect 391 151 393 156
rect 401 151 403 156
rect 439 164 441 173
rect 461 164 463 173
rect 472 170 474 173
rect 479 170 481 173
rect 499 170 501 173
rect 509 170 511 173
rect 519 178 521 180
rect 523 178 525 180
rect 519 176 525 178
rect 519 163 521 176
rect 529 172 531 185
rect 546 184 552 186
rect 546 182 548 184
rect 550 182 552 184
rect 546 180 552 182
rect 525 170 531 172
rect 550 170 552 180
rect 557 179 559 189
rect 618 201 620 205
rect 598 187 600 190
rect 594 185 600 187
rect 594 183 596 185
rect 598 183 600 185
rect 570 179 572 182
rect 594 181 600 183
rect 556 177 562 179
rect 556 175 558 177
rect 560 175 562 177
rect 556 173 562 175
rect 566 177 572 179
rect 566 175 568 177
rect 570 175 572 177
rect 566 173 572 175
rect 560 170 562 173
rect 570 170 572 173
rect 525 168 527 170
rect 529 168 531 170
rect 525 166 531 168
rect 529 163 531 166
rect 499 151 501 156
rect 509 151 511 156
rect 421 146 423 150
rect 428 146 430 150
rect 439 146 441 150
rect 461 146 463 150
rect 472 146 474 150
rect 479 146 481 150
rect 519 148 521 153
rect 550 159 552 164
rect 560 159 562 164
rect 598 168 600 181
rect 608 179 610 190
rect 670 207 672 212
rect 677 207 679 212
rect 695 210 697 214
rect 705 210 707 214
rect 715 210 717 214
rect 737 210 739 214
rect 747 210 749 214
rect 757 210 759 214
rect 660 198 662 203
rect 618 179 620 183
rect 604 177 610 179
rect 604 175 606 177
rect 608 175 610 177
rect 604 173 610 175
rect 614 177 620 179
rect 614 175 616 177
rect 618 175 620 177
rect 614 173 620 175
rect 605 168 607 173
rect 618 168 620 173
rect 647 172 649 185
rect 660 182 662 185
rect 775 207 777 212
rect 782 207 784 212
rect 805 210 807 214
rect 826 210 828 214
rect 833 210 835 214
rect 792 198 794 203
rect 924 210 926 214
rect 846 200 848 205
rect 874 203 876 208
rect 884 203 886 208
rect 826 186 828 189
rect 792 182 794 185
rect 653 180 662 182
rect 653 178 655 180
rect 657 178 659 180
rect 670 179 672 182
rect 677 179 679 182
rect 695 179 697 182
rect 705 179 707 182
rect 715 179 717 182
rect 737 179 739 182
rect 747 179 749 182
rect 757 179 759 182
rect 775 179 777 182
rect 782 179 784 182
rect 792 180 801 182
rect 653 176 659 178
rect 647 170 653 172
rect 647 168 649 170
rect 651 168 653 170
rect 570 156 572 161
rect 647 166 653 168
rect 647 163 649 166
rect 657 163 659 176
rect 667 177 673 179
rect 667 175 669 177
rect 671 175 673 177
rect 667 173 673 175
rect 677 177 699 179
rect 677 175 688 177
rect 690 175 695 177
rect 697 175 699 177
rect 677 173 699 175
rect 703 177 709 179
rect 703 175 705 177
rect 707 175 709 177
rect 703 173 709 175
rect 713 177 719 179
rect 713 175 715 177
rect 717 175 719 177
rect 713 173 719 175
rect 735 177 741 179
rect 735 175 737 177
rect 739 175 741 177
rect 735 173 741 175
rect 745 177 751 179
rect 745 175 747 177
rect 749 175 751 177
rect 745 173 751 175
rect 755 177 777 179
rect 755 175 757 177
rect 759 175 764 177
rect 766 175 777 177
rect 755 173 777 175
rect 781 177 787 179
rect 781 175 783 177
rect 785 175 787 177
rect 781 173 787 175
rect 667 170 669 173
rect 677 170 679 173
rect 697 170 699 173
rect 704 170 706 173
rect 598 152 600 157
rect 605 152 607 157
rect 529 146 531 150
rect 618 155 620 159
rect 647 146 649 150
rect 657 148 659 153
rect 667 151 669 156
rect 677 151 679 156
rect 715 164 717 173
rect 737 164 739 173
rect 748 170 750 173
rect 755 170 757 173
rect 775 170 777 173
rect 785 170 787 173
rect 795 178 797 180
rect 799 178 801 180
rect 795 176 801 178
rect 795 163 797 176
rect 805 172 807 185
rect 822 184 828 186
rect 822 182 824 184
rect 826 182 828 184
rect 822 180 828 182
rect 801 170 807 172
rect 826 170 828 180
rect 833 179 835 189
rect 894 201 896 205
rect 874 187 876 190
rect 870 185 876 187
rect 870 183 872 185
rect 874 183 876 185
rect 846 179 848 182
rect 870 181 876 183
rect 832 177 838 179
rect 832 175 834 177
rect 836 175 838 177
rect 832 173 838 175
rect 842 177 848 179
rect 842 175 844 177
rect 846 175 848 177
rect 842 173 848 175
rect 836 170 838 173
rect 846 170 848 173
rect 801 168 803 170
rect 805 168 807 170
rect 801 166 807 168
rect 805 163 807 166
rect 775 151 777 156
rect 785 151 787 156
rect 697 146 699 150
rect 704 146 706 150
rect 715 146 717 150
rect 737 146 739 150
rect 748 146 750 150
rect 755 146 757 150
rect 795 148 797 153
rect 826 159 828 164
rect 836 159 838 164
rect 874 168 876 181
rect 884 179 886 190
rect 947 207 949 212
rect 954 207 956 212
rect 972 210 974 214
rect 982 210 984 214
rect 992 210 994 214
rect 1014 210 1016 214
rect 1024 210 1026 214
rect 1034 210 1036 214
rect 937 198 939 203
rect 894 179 896 183
rect 880 177 886 179
rect 880 175 882 177
rect 884 175 886 177
rect 880 173 886 175
rect 890 177 896 179
rect 890 175 892 177
rect 894 175 896 177
rect 890 173 896 175
rect 881 168 883 173
rect 894 168 896 173
rect 924 172 926 185
rect 937 182 939 185
rect 1052 207 1054 212
rect 1059 207 1061 212
rect 1082 210 1084 214
rect 1103 210 1105 214
rect 1110 210 1112 214
rect 1069 198 1071 203
rect 1123 200 1125 205
rect 1103 186 1105 189
rect 1069 182 1071 185
rect 930 180 939 182
rect 930 178 932 180
rect 934 178 936 180
rect 947 179 949 182
rect 954 179 956 182
rect 972 179 974 182
rect 982 179 984 182
rect 992 179 994 182
rect 1014 179 1016 182
rect 1024 179 1026 182
rect 1034 179 1036 182
rect 1052 179 1054 182
rect 1059 179 1061 182
rect 1069 180 1078 182
rect 930 176 936 178
rect 924 170 930 172
rect 924 168 926 170
rect 928 168 930 170
rect 846 156 848 161
rect 924 166 930 168
rect 924 163 926 166
rect 934 163 936 176
rect 944 177 950 179
rect 944 175 946 177
rect 948 175 950 177
rect 944 173 950 175
rect 954 177 976 179
rect 954 175 965 177
rect 967 175 972 177
rect 974 175 976 177
rect 954 173 976 175
rect 980 177 986 179
rect 980 175 982 177
rect 984 175 986 177
rect 980 173 986 175
rect 990 177 996 179
rect 990 175 992 177
rect 994 175 996 177
rect 990 173 996 175
rect 1012 177 1018 179
rect 1012 175 1014 177
rect 1016 175 1018 177
rect 1012 173 1018 175
rect 1022 177 1028 179
rect 1022 175 1024 177
rect 1026 175 1028 177
rect 1022 173 1028 175
rect 1032 177 1054 179
rect 1032 175 1034 177
rect 1036 175 1041 177
rect 1043 175 1054 177
rect 1032 173 1054 175
rect 1058 177 1064 179
rect 1058 175 1060 177
rect 1062 175 1064 177
rect 1058 173 1064 175
rect 944 170 946 173
rect 954 170 956 173
rect 974 170 976 173
rect 981 170 983 173
rect 874 152 876 157
rect 881 152 883 157
rect 805 146 807 150
rect 894 155 896 159
rect 924 146 926 150
rect 934 148 936 153
rect 944 151 946 156
rect 954 151 956 156
rect 992 164 994 173
rect 1014 164 1016 173
rect 1025 170 1027 173
rect 1032 170 1034 173
rect 1052 170 1054 173
rect 1062 170 1064 173
rect 1072 178 1074 180
rect 1076 178 1078 180
rect 1072 176 1078 178
rect 1072 163 1074 176
rect 1082 172 1084 185
rect 1099 184 1105 186
rect 1099 182 1101 184
rect 1103 182 1105 184
rect 1099 180 1105 182
rect 1078 170 1084 172
rect 1103 170 1105 180
rect 1110 179 1112 189
rect 1123 179 1125 182
rect 1109 177 1115 179
rect 1109 175 1111 177
rect 1113 175 1115 177
rect 1109 173 1115 175
rect 1119 177 1125 179
rect 1119 175 1121 177
rect 1123 175 1125 177
rect 1119 173 1125 175
rect 1113 170 1115 173
rect 1123 170 1125 173
rect 1078 168 1080 170
rect 1082 168 1084 170
rect 1078 166 1084 168
rect 1082 163 1084 166
rect 1052 151 1054 156
rect 1062 151 1064 156
rect 974 146 976 150
rect 981 146 983 150
rect 992 146 994 150
rect 1014 146 1016 150
rect 1025 146 1027 150
rect 1032 146 1034 150
rect 1072 148 1074 153
rect 1103 159 1105 164
rect 1113 159 1115 164
rect 1123 156 1125 161
rect 1082 146 1084 150
rect -273 140 -248 142
rect -273 132 -271 140
rect -260 132 -258 136
rect -250 132 -248 140
rect -240 135 -238 140
rect -233 135 -231 140
rect -208 138 -206 142
rect -276 130 -271 132
rect -276 127 -274 130
rect -198 135 -196 140
rect -158 138 -156 142
rect -151 138 -149 142
rect -140 138 -138 142
rect -118 138 -116 142
rect -107 138 -105 142
rect -100 138 -98 142
rect -188 132 -186 137
rect -178 132 -176 137
rect -260 120 -258 123
rect -267 118 -258 120
rect -250 119 -248 123
rect -240 120 -238 123
rect -276 110 -274 118
rect -267 116 -265 118
rect -263 116 -258 118
rect -267 114 -258 116
rect -242 118 -238 120
rect -242 115 -240 118
rect -260 110 -258 114
rect -246 113 -240 115
rect -233 114 -231 123
rect -208 122 -206 125
rect -208 120 -202 122
rect -208 118 -206 120
rect -204 118 -202 120
rect -208 116 -202 118
rect -246 111 -244 113
rect -242 111 -240 113
rect -279 108 -266 110
rect -260 108 -250 110
rect -246 109 -240 111
rect -279 107 -277 108
rect -283 105 -277 107
rect -268 105 -266 108
rect -252 105 -250 108
rect -242 105 -240 109
rect -236 112 -230 114
rect -236 110 -234 112
rect -232 110 -230 112
rect -236 108 -230 110
rect -232 105 -230 108
rect -283 103 -281 105
rect -279 103 -277 105
rect -283 101 -277 103
rect -252 83 -250 87
rect -242 83 -240 87
rect -268 74 -266 78
rect -208 103 -206 116
rect -198 112 -196 125
rect -202 110 -196 112
rect -202 108 -200 110
rect -198 108 -196 110
rect -188 115 -186 118
rect -178 115 -176 118
rect -158 115 -156 118
rect -151 115 -149 118
rect -140 115 -138 124
rect -118 115 -116 124
rect -80 132 -78 137
rect -70 132 -68 137
rect -60 135 -58 140
rect -50 138 -48 142
rect -107 115 -105 118
rect -100 115 -98 118
rect -80 115 -78 118
rect -70 115 -68 118
rect -188 113 -182 115
rect -188 111 -186 113
rect -184 111 -182 113
rect -188 109 -182 111
rect -178 113 -156 115
rect -178 111 -167 113
rect -165 111 -160 113
rect -158 111 -156 113
rect -178 109 -156 111
rect -152 113 -146 115
rect -152 111 -150 113
rect -148 111 -146 113
rect -152 109 -146 111
rect -142 113 -136 115
rect -142 111 -140 113
rect -138 111 -136 113
rect -142 109 -136 111
rect -120 113 -114 115
rect -120 111 -118 113
rect -116 111 -114 113
rect -120 109 -114 111
rect -110 113 -104 115
rect -110 111 -108 113
rect -106 111 -104 113
rect -110 109 -104 111
rect -100 113 -78 115
rect -100 111 -98 113
rect -96 111 -91 113
rect -89 111 -78 113
rect -100 109 -78 111
rect -74 113 -68 115
rect -74 111 -72 113
rect -70 111 -68 113
rect -74 109 -68 111
rect -60 112 -58 125
rect -50 122 -48 125
rect -54 120 -48 122
rect -54 118 -52 120
rect -50 118 -48 120
rect -29 124 -27 129
rect -19 124 -17 129
rect -9 127 -7 132
rect 14 131 16 136
rect 21 131 23 136
rect 34 129 36 133
rect 54 131 56 136
rect 61 131 63 136
rect 94 138 96 142
rect 74 129 76 133
rect 104 135 106 140
rect 144 138 146 142
rect 151 138 153 142
rect 162 138 164 142
rect 184 138 186 142
rect 195 138 197 142
rect 202 138 204 142
rect 114 132 116 137
rect 124 132 126 137
rect 94 122 96 125
rect 94 120 100 122
rect -54 116 -48 118
rect -60 110 -54 112
rect -202 106 -193 108
rect -185 106 -183 109
rect -178 106 -176 109
rect -160 106 -158 109
rect -150 106 -148 109
rect -140 106 -138 109
rect -118 106 -116 109
rect -108 106 -106 109
rect -98 106 -96 109
rect -80 106 -78 109
rect -73 106 -71 109
rect -60 108 -58 110
rect -56 108 -54 110
rect -63 106 -54 108
rect -195 103 -193 106
rect -195 85 -193 90
rect -232 74 -230 78
rect -208 74 -206 78
rect -185 76 -183 81
rect -178 76 -176 81
rect -63 103 -61 106
rect -50 103 -48 116
rect -29 108 -27 118
rect -19 115 -17 118
rect -9 115 -7 118
rect -23 113 -17 115
rect -23 111 -21 113
rect -19 111 -17 113
rect -23 109 -17 111
rect -13 113 -7 115
rect -13 111 -11 113
rect -9 111 -7 113
rect -13 109 -7 111
rect -33 106 -27 108
rect -33 104 -31 106
rect -29 104 -27 106
rect -63 85 -61 90
rect -160 74 -158 78
rect -150 74 -148 78
rect -140 74 -138 78
rect -118 74 -116 78
rect -108 74 -106 78
rect -98 74 -96 78
rect -80 76 -78 81
rect -73 76 -71 81
rect -33 102 -27 104
rect -29 99 -27 102
rect -22 99 -20 109
rect -9 106 -7 109
rect 14 107 16 120
rect 21 115 23 120
rect 34 115 36 120
rect 20 113 26 115
rect 20 111 22 113
rect 24 111 26 113
rect 20 109 26 111
rect 30 113 36 115
rect 30 111 32 113
rect 34 111 36 113
rect 30 109 36 111
rect 10 105 16 107
rect 10 103 12 105
rect 14 103 16 105
rect 10 101 16 103
rect 14 98 16 101
rect 24 98 26 109
rect 34 105 36 109
rect 54 107 56 120
rect 61 115 63 120
rect 74 115 76 120
rect 60 113 66 115
rect 60 111 62 113
rect 64 111 66 113
rect 60 109 66 111
rect 70 113 76 115
rect 70 111 72 113
rect 74 111 76 113
rect 70 109 76 111
rect 50 105 56 107
rect -9 83 -7 88
rect 50 103 52 105
rect 54 103 56 105
rect 50 101 56 103
rect 54 98 56 101
rect 64 98 66 109
rect 74 105 76 109
rect 94 118 96 120
rect 98 118 100 120
rect 94 116 100 118
rect 14 80 16 85
rect 24 80 26 85
rect 34 83 36 87
rect 94 103 96 116
rect 104 112 106 125
rect 100 110 106 112
rect 100 108 102 110
rect 104 108 106 110
rect 114 115 116 118
rect 124 115 126 118
rect 144 115 146 118
rect 151 115 153 118
rect 162 115 164 124
rect 184 115 186 124
rect 222 132 224 137
rect 232 132 234 137
rect 242 135 244 140
rect 252 138 254 142
rect 195 115 197 118
rect 202 115 204 118
rect 222 115 224 118
rect 232 115 234 118
rect 114 113 120 115
rect 114 111 116 113
rect 118 111 120 113
rect 114 109 120 111
rect 124 113 146 115
rect 124 111 135 113
rect 137 111 142 113
rect 144 111 146 113
rect 124 109 146 111
rect 150 113 156 115
rect 150 111 152 113
rect 154 111 156 113
rect 150 109 156 111
rect 160 113 166 115
rect 160 111 162 113
rect 164 111 166 113
rect 160 109 166 111
rect 182 113 188 115
rect 182 111 184 113
rect 186 111 188 113
rect 182 109 188 111
rect 192 113 198 115
rect 192 111 194 113
rect 196 111 198 113
rect 192 109 198 111
rect 202 113 224 115
rect 202 111 204 113
rect 206 111 211 113
rect 213 111 224 113
rect 202 109 224 111
rect 228 113 234 115
rect 228 111 230 113
rect 232 111 234 113
rect 228 109 234 111
rect 242 112 244 125
rect 252 122 254 125
rect 248 120 254 122
rect 248 118 250 120
rect 252 118 254 120
rect 273 124 275 129
rect 283 124 285 129
rect 293 127 295 132
rect 321 131 323 136
rect 328 131 330 136
rect 371 138 373 142
rect 341 129 343 133
rect 381 135 383 140
rect 421 138 423 142
rect 428 138 430 142
rect 439 138 441 142
rect 461 138 463 142
rect 472 138 474 142
rect 479 138 481 142
rect 391 132 393 137
rect 401 132 403 137
rect 371 122 373 125
rect 371 120 377 122
rect 248 116 254 118
rect 242 110 248 112
rect 100 106 109 108
rect 117 106 119 109
rect 124 106 126 109
rect 142 106 144 109
rect 152 106 154 109
rect 162 106 164 109
rect 184 106 186 109
rect 194 106 196 109
rect 204 106 206 109
rect 222 106 224 109
rect 229 106 231 109
rect 242 108 244 110
rect 246 108 248 110
rect 239 106 248 108
rect 107 103 109 106
rect -50 74 -48 78
rect -29 74 -27 78
rect -22 74 -20 78
rect 54 80 56 85
rect 64 80 66 85
rect 74 83 76 87
rect 107 85 109 90
rect 94 74 96 78
rect 117 76 119 81
rect 124 76 126 81
rect 239 103 241 106
rect 252 103 254 116
rect 273 108 275 118
rect 283 115 285 118
rect 293 115 295 118
rect 279 113 285 115
rect 279 111 281 113
rect 283 111 285 113
rect 279 109 285 111
rect 289 113 295 115
rect 289 111 291 113
rect 293 111 295 113
rect 289 109 295 111
rect 269 106 275 108
rect 269 104 271 106
rect 273 104 275 106
rect 239 85 241 90
rect 142 74 144 78
rect 152 74 154 78
rect 162 74 164 78
rect 184 74 186 78
rect 194 74 196 78
rect 204 74 206 78
rect 222 76 224 81
rect 229 76 231 81
rect 269 102 275 104
rect 273 99 275 102
rect 280 99 282 109
rect 293 106 295 109
rect 321 107 323 120
rect 328 115 330 120
rect 341 115 343 120
rect 327 113 333 115
rect 327 111 329 113
rect 331 111 333 113
rect 327 109 333 111
rect 337 113 343 115
rect 337 111 339 113
rect 341 111 343 113
rect 337 109 343 111
rect 317 105 323 107
rect 317 103 319 105
rect 321 103 323 105
rect 317 101 323 103
rect 321 98 323 101
rect 331 98 333 109
rect 341 105 343 109
rect 371 118 373 120
rect 375 118 377 120
rect 371 116 377 118
rect 293 83 295 88
rect 371 103 373 116
rect 381 112 383 125
rect 377 110 383 112
rect 377 108 379 110
rect 381 108 383 110
rect 391 115 393 118
rect 401 115 403 118
rect 421 115 423 118
rect 428 115 430 118
rect 439 115 441 124
rect 461 115 463 124
rect 499 132 501 137
rect 509 132 511 137
rect 519 135 521 140
rect 529 138 531 142
rect 472 115 474 118
rect 479 115 481 118
rect 499 115 501 118
rect 509 115 511 118
rect 391 113 397 115
rect 391 111 393 113
rect 395 111 397 113
rect 391 109 397 111
rect 401 113 423 115
rect 401 111 412 113
rect 414 111 419 113
rect 421 111 423 113
rect 401 109 423 111
rect 427 113 433 115
rect 427 111 429 113
rect 431 111 433 113
rect 427 109 433 111
rect 437 113 443 115
rect 437 111 439 113
rect 441 111 443 113
rect 437 109 443 111
rect 459 113 465 115
rect 459 111 461 113
rect 463 111 465 113
rect 459 109 465 111
rect 469 113 475 115
rect 469 111 471 113
rect 473 111 475 113
rect 469 109 475 111
rect 479 113 501 115
rect 479 111 481 113
rect 483 111 488 113
rect 490 111 501 113
rect 479 109 501 111
rect 505 113 511 115
rect 505 111 507 113
rect 509 111 511 113
rect 505 109 511 111
rect 519 112 521 125
rect 529 122 531 125
rect 525 120 531 122
rect 525 118 527 120
rect 529 118 531 120
rect 550 124 552 129
rect 560 124 562 129
rect 570 127 572 132
rect 598 131 600 136
rect 605 131 607 136
rect 647 138 649 142
rect 618 129 620 133
rect 657 135 659 140
rect 697 138 699 142
rect 704 138 706 142
rect 715 138 717 142
rect 737 138 739 142
rect 748 138 750 142
rect 755 138 757 142
rect 667 132 669 137
rect 677 132 679 137
rect 647 122 649 125
rect 647 120 653 122
rect 525 116 531 118
rect 519 110 525 112
rect 377 106 386 108
rect 394 106 396 109
rect 401 106 403 109
rect 419 106 421 109
rect 429 106 431 109
rect 439 106 441 109
rect 461 106 463 109
rect 471 106 473 109
rect 481 106 483 109
rect 499 106 501 109
rect 506 106 508 109
rect 519 108 521 110
rect 523 108 525 110
rect 516 106 525 108
rect 384 103 386 106
rect 321 80 323 85
rect 331 80 333 85
rect 341 83 343 87
rect 252 74 254 78
rect 273 74 275 78
rect 280 74 282 78
rect 384 85 386 90
rect 371 74 373 78
rect 394 76 396 81
rect 401 76 403 81
rect 516 103 518 106
rect 529 103 531 116
rect 550 108 552 118
rect 560 115 562 118
rect 570 115 572 118
rect 556 113 562 115
rect 556 111 558 113
rect 560 111 562 113
rect 556 109 562 111
rect 566 113 572 115
rect 566 111 568 113
rect 570 111 572 113
rect 566 109 572 111
rect 546 106 552 108
rect 546 104 548 106
rect 550 104 552 106
rect 516 85 518 90
rect 419 74 421 78
rect 429 74 431 78
rect 439 74 441 78
rect 461 74 463 78
rect 471 74 473 78
rect 481 74 483 78
rect 499 76 501 81
rect 506 76 508 81
rect 546 102 552 104
rect 550 99 552 102
rect 557 99 559 109
rect 570 106 572 109
rect 598 107 600 120
rect 605 115 607 120
rect 618 115 620 120
rect 604 113 610 115
rect 604 111 606 113
rect 608 111 610 113
rect 604 109 610 111
rect 614 113 620 115
rect 614 111 616 113
rect 618 111 620 113
rect 614 109 620 111
rect 594 105 600 107
rect 594 103 596 105
rect 598 103 600 105
rect 594 101 600 103
rect 598 98 600 101
rect 608 98 610 109
rect 618 105 620 109
rect 647 118 649 120
rect 651 118 653 120
rect 647 116 653 118
rect 570 83 572 88
rect 647 103 649 116
rect 657 112 659 125
rect 653 110 659 112
rect 653 108 655 110
rect 657 108 659 110
rect 667 115 669 118
rect 677 115 679 118
rect 697 115 699 118
rect 704 115 706 118
rect 715 115 717 124
rect 737 115 739 124
rect 775 132 777 137
rect 785 132 787 137
rect 795 135 797 140
rect 805 138 807 142
rect 748 115 750 118
rect 755 115 757 118
rect 775 115 777 118
rect 785 115 787 118
rect 667 113 673 115
rect 667 111 669 113
rect 671 111 673 113
rect 667 109 673 111
rect 677 113 699 115
rect 677 111 688 113
rect 690 111 695 113
rect 697 111 699 113
rect 677 109 699 111
rect 703 113 709 115
rect 703 111 705 113
rect 707 111 709 113
rect 703 109 709 111
rect 713 113 719 115
rect 713 111 715 113
rect 717 111 719 113
rect 713 109 719 111
rect 735 113 741 115
rect 735 111 737 113
rect 739 111 741 113
rect 735 109 741 111
rect 745 113 751 115
rect 745 111 747 113
rect 749 111 751 113
rect 745 109 751 111
rect 755 113 777 115
rect 755 111 757 113
rect 759 111 764 113
rect 766 111 777 113
rect 755 109 777 111
rect 781 113 787 115
rect 781 111 783 113
rect 785 111 787 113
rect 781 109 787 111
rect 795 112 797 125
rect 805 122 807 125
rect 801 120 807 122
rect 801 118 803 120
rect 805 118 807 120
rect 826 124 828 129
rect 836 124 838 129
rect 846 127 848 132
rect 874 131 876 136
rect 881 131 883 136
rect 924 138 926 142
rect 894 129 896 133
rect 934 135 936 140
rect 974 138 976 142
rect 981 138 983 142
rect 992 138 994 142
rect 1014 138 1016 142
rect 1025 138 1027 142
rect 1032 138 1034 142
rect 944 132 946 137
rect 954 132 956 137
rect 924 122 926 125
rect 924 120 930 122
rect 801 116 807 118
rect 795 110 801 112
rect 653 106 662 108
rect 670 106 672 109
rect 677 106 679 109
rect 695 106 697 109
rect 705 106 707 109
rect 715 106 717 109
rect 737 106 739 109
rect 747 106 749 109
rect 757 106 759 109
rect 775 106 777 109
rect 782 106 784 109
rect 795 108 797 110
rect 799 108 801 110
rect 792 106 801 108
rect 660 103 662 106
rect 598 80 600 85
rect 608 80 610 85
rect 618 83 620 87
rect 529 74 531 78
rect 550 74 552 78
rect 557 74 559 78
rect 660 85 662 90
rect 647 74 649 78
rect 670 76 672 81
rect 677 76 679 81
rect 792 103 794 106
rect 805 103 807 116
rect 826 108 828 118
rect 836 115 838 118
rect 846 115 848 118
rect 832 113 838 115
rect 832 111 834 113
rect 836 111 838 113
rect 832 109 838 111
rect 842 113 848 115
rect 842 111 844 113
rect 846 111 848 113
rect 842 109 848 111
rect 822 106 828 108
rect 822 104 824 106
rect 826 104 828 106
rect 792 85 794 90
rect 695 74 697 78
rect 705 74 707 78
rect 715 74 717 78
rect 737 74 739 78
rect 747 74 749 78
rect 757 74 759 78
rect 775 76 777 81
rect 782 76 784 81
rect 822 102 828 104
rect 826 99 828 102
rect 833 99 835 109
rect 846 106 848 109
rect 874 107 876 120
rect 881 115 883 120
rect 894 115 896 120
rect 880 113 886 115
rect 880 111 882 113
rect 884 111 886 113
rect 880 109 886 111
rect 890 113 896 115
rect 890 111 892 113
rect 894 111 896 113
rect 890 109 896 111
rect 870 105 876 107
rect 870 103 872 105
rect 874 103 876 105
rect 870 101 876 103
rect 874 98 876 101
rect 884 98 886 109
rect 894 105 896 109
rect 924 118 926 120
rect 928 118 930 120
rect 924 116 930 118
rect 846 83 848 88
rect 924 103 926 116
rect 934 112 936 125
rect 930 110 936 112
rect 930 108 932 110
rect 934 108 936 110
rect 944 115 946 118
rect 954 115 956 118
rect 974 115 976 118
rect 981 115 983 118
rect 992 115 994 124
rect 1014 115 1016 124
rect 1052 132 1054 137
rect 1062 132 1064 137
rect 1072 135 1074 140
rect 1082 138 1084 142
rect 1025 115 1027 118
rect 1032 115 1034 118
rect 1052 115 1054 118
rect 1062 115 1064 118
rect 944 113 950 115
rect 944 111 946 113
rect 948 111 950 113
rect 944 109 950 111
rect 954 113 976 115
rect 954 111 965 113
rect 967 111 972 113
rect 974 111 976 113
rect 954 109 976 111
rect 980 113 986 115
rect 980 111 982 113
rect 984 111 986 113
rect 980 109 986 111
rect 990 113 996 115
rect 990 111 992 113
rect 994 111 996 113
rect 990 109 996 111
rect 1012 113 1018 115
rect 1012 111 1014 113
rect 1016 111 1018 113
rect 1012 109 1018 111
rect 1022 113 1028 115
rect 1022 111 1024 113
rect 1026 111 1028 113
rect 1022 109 1028 111
rect 1032 113 1054 115
rect 1032 111 1034 113
rect 1036 111 1041 113
rect 1043 111 1054 113
rect 1032 109 1054 111
rect 1058 113 1064 115
rect 1058 111 1060 113
rect 1062 111 1064 113
rect 1058 109 1064 111
rect 1072 112 1074 125
rect 1082 122 1084 125
rect 1078 120 1084 122
rect 1078 118 1080 120
rect 1082 118 1084 120
rect 1103 124 1105 129
rect 1113 124 1115 129
rect 1123 127 1125 132
rect 1078 116 1084 118
rect 1072 110 1078 112
rect 930 106 939 108
rect 947 106 949 109
rect 954 106 956 109
rect 972 106 974 109
rect 982 106 984 109
rect 992 106 994 109
rect 1014 106 1016 109
rect 1024 106 1026 109
rect 1034 106 1036 109
rect 1052 106 1054 109
rect 1059 106 1061 109
rect 1072 108 1074 110
rect 1076 108 1078 110
rect 1069 106 1078 108
rect 937 103 939 106
rect 874 80 876 85
rect 884 80 886 85
rect 894 83 896 87
rect 805 74 807 78
rect 826 74 828 78
rect 833 74 835 78
rect 937 85 939 90
rect 924 74 926 78
rect 947 76 949 81
rect 954 76 956 81
rect 1069 103 1071 106
rect 1082 103 1084 116
rect 1103 108 1105 118
rect 1113 115 1115 118
rect 1123 115 1125 118
rect 1109 113 1115 115
rect 1109 111 1111 113
rect 1113 111 1115 113
rect 1109 109 1115 111
rect 1119 113 1125 115
rect 1119 111 1121 113
rect 1123 111 1125 113
rect 1119 109 1125 111
rect 1099 106 1105 108
rect 1099 104 1101 106
rect 1103 104 1105 106
rect 1069 85 1071 90
rect 972 74 974 78
rect 982 74 984 78
rect 992 74 994 78
rect 1014 74 1016 78
rect 1024 74 1026 78
rect 1034 74 1036 78
rect 1052 76 1054 81
rect 1059 76 1061 81
rect 1099 102 1105 104
rect 1103 99 1105 102
rect 1110 99 1112 109
rect 1123 106 1125 109
rect 1123 83 1125 88
rect 1082 74 1084 78
rect 1103 74 1105 78
rect 1110 74 1112 78
rect -268 66 -266 70
rect -283 41 -277 43
rect -283 39 -281 41
rect -279 39 -277 41
rect -232 66 -230 70
rect -208 66 -206 70
rect -252 57 -250 61
rect -242 57 -240 61
rect -185 63 -183 68
rect -178 63 -176 68
rect -160 66 -158 70
rect -150 66 -148 70
rect -140 66 -138 70
rect -118 66 -116 70
rect -108 66 -106 70
rect -98 66 -96 70
rect -195 54 -193 59
rect -283 37 -277 39
rect -279 36 -277 37
rect -268 36 -266 39
rect -252 36 -250 39
rect -279 34 -266 36
rect -260 34 -250 36
rect -242 35 -240 39
rect -232 36 -230 39
rect -276 26 -274 34
rect -260 30 -258 34
rect -267 28 -258 30
rect -246 33 -240 35
rect -246 31 -244 33
rect -242 31 -240 33
rect -246 29 -240 31
rect -236 34 -230 36
rect -236 32 -234 34
rect -232 32 -230 34
rect -236 30 -230 32
rect -267 26 -265 28
rect -263 26 -258 28
rect -267 24 -258 26
rect -242 26 -240 29
rect -260 21 -258 24
rect -250 21 -248 25
rect -242 24 -238 26
rect -240 21 -238 24
rect -233 21 -231 30
rect -208 28 -206 41
rect -195 38 -193 41
rect -80 63 -78 68
rect -73 63 -71 68
rect -50 66 -48 70
rect -29 66 -27 70
rect -22 66 -20 70
rect -63 54 -61 59
rect -9 56 -7 61
rect 14 59 16 64
rect 24 59 26 64
rect 94 66 96 70
rect -29 42 -27 45
rect -63 38 -61 41
rect -202 36 -193 38
rect -202 34 -200 36
rect -198 34 -196 36
rect -185 35 -183 38
rect -178 35 -176 38
rect -160 35 -158 38
rect -150 35 -148 38
rect -140 35 -138 38
rect -118 35 -116 38
rect -108 35 -106 38
rect -98 35 -96 38
rect -80 35 -78 38
rect -73 35 -71 38
rect -63 36 -54 38
rect -202 32 -196 34
rect -208 26 -202 28
rect -208 24 -206 26
rect -204 24 -202 26
rect -208 22 -202 24
rect -276 14 -274 17
rect -276 12 -271 14
rect -273 4 -271 12
rect -260 8 -258 12
rect -250 4 -248 12
rect -208 19 -206 22
rect -198 19 -196 32
rect -188 33 -182 35
rect -188 31 -186 33
rect -184 31 -182 33
rect -188 29 -182 31
rect -178 33 -156 35
rect -178 31 -167 33
rect -165 31 -160 33
rect -158 31 -156 33
rect -178 29 -156 31
rect -152 33 -146 35
rect -152 31 -150 33
rect -148 31 -146 33
rect -152 29 -146 31
rect -142 33 -136 35
rect -142 31 -140 33
rect -138 31 -136 33
rect -142 29 -136 31
rect -120 33 -114 35
rect -120 31 -118 33
rect -116 31 -114 33
rect -120 29 -114 31
rect -110 33 -104 35
rect -110 31 -108 33
rect -106 31 -104 33
rect -110 29 -104 31
rect -100 33 -78 35
rect -100 31 -98 33
rect -96 31 -91 33
rect -89 31 -78 33
rect -100 29 -78 31
rect -74 33 -68 35
rect -74 31 -72 33
rect -70 31 -68 33
rect -74 29 -68 31
rect -188 26 -186 29
rect -178 26 -176 29
rect -158 26 -156 29
rect -151 26 -149 29
rect -240 4 -238 9
rect -233 4 -231 9
rect -273 2 -248 4
rect -208 2 -206 6
rect -198 4 -196 9
rect -188 7 -186 12
rect -178 7 -176 12
rect -140 20 -138 29
rect -118 20 -116 29
rect -107 26 -105 29
rect -100 26 -98 29
rect -80 26 -78 29
rect -70 26 -68 29
rect -60 34 -58 36
rect -56 34 -54 36
rect -60 32 -54 34
rect -60 19 -58 32
rect -50 28 -48 41
rect -33 40 -27 42
rect -33 38 -31 40
rect -29 38 -27 40
rect -33 36 -27 38
rect -54 26 -48 28
rect -29 26 -27 36
rect -22 35 -20 45
rect 34 57 36 61
rect 54 59 56 64
rect 64 59 66 64
rect 14 43 16 46
rect 10 41 16 43
rect 10 39 12 41
rect 14 39 16 41
rect -9 35 -7 38
rect 10 37 16 39
rect -23 33 -17 35
rect -23 31 -21 33
rect -19 31 -17 33
rect -23 29 -17 31
rect -13 33 -7 35
rect -13 31 -11 33
rect -9 31 -7 33
rect -13 29 -7 31
rect -19 26 -17 29
rect -9 26 -7 29
rect -54 24 -52 26
rect -50 24 -48 26
rect -54 22 -48 24
rect -50 19 -48 22
rect -80 7 -78 12
rect -70 7 -68 12
rect -158 2 -156 6
rect -151 2 -149 6
rect -140 2 -138 6
rect -118 2 -116 6
rect -107 2 -105 6
rect -100 2 -98 6
rect -60 4 -58 9
rect -29 15 -27 20
rect -19 15 -17 20
rect 14 24 16 37
rect 24 35 26 46
rect 74 57 76 61
rect 54 43 56 46
rect 50 41 56 43
rect 50 39 52 41
rect 54 39 56 41
rect 34 35 36 39
rect 50 37 56 39
rect 20 33 26 35
rect 20 31 22 33
rect 24 31 26 33
rect 20 29 26 31
rect 30 33 36 35
rect 30 31 32 33
rect 34 31 36 33
rect 30 29 36 31
rect 21 24 23 29
rect 34 24 36 29
rect 54 24 56 37
rect 64 35 66 46
rect 117 63 119 68
rect 124 63 126 68
rect 142 66 144 70
rect 152 66 154 70
rect 162 66 164 70
rect 184 66 186 70
rect 194 66 196 70
rect 204 66 206 70
rect 107 54 109 59
rect 74 35 76 39
rect 60 33 66 35
rect 60 31 62 33
rect 64 31 66 33
rect 60 29 66 31
rect 70 33 76 35
rect 70 31 72 33
rect 74 31 76 33
rect 70 29 76 31
rect 61 24 63 29
rect 74 24 76 29
rect 94 28 96 41
rect 107 38 109 41
rect 222 63 224 68
rect 229 63 231 68
rect 252 66 254 70
rect 273 66 275 70
rect 280 66 282 70
rect 239 54 241 59
rect 371 66 373 70
rect 293 56 295 61
rect 321 59 323 64
rect 331 59 333 64
rect 273 42 275 45
rect 239 38 241 41
rect 100 36 109 38
rect 100 34 102 36
rect 104 34 106 36
rect 117 35 119 38
rect 124 35 126 38
rect 142 35 144 38
rect 152 35 154 38
rect 162 35 164 38
rect 184 35 186 38
rect 194 35 196 38
rect 204 35 206 38
rect 222 35 224 38
rect 229 35 231 38
rect 239 36 248 38
rect 100 32 106 34
rect 94 26 100 28
rect 94 24 96 26
rect 98 24 100 26
rect -9 12 -7 17
rect 14 8 16 13
rect 21 8 23 13
rect -50 2 -48 6
rect 34 11 36 15
rect 94 22 100 24
rect 94 19 96 22
rect 104 19 106 32
rect 114 33 120 35
rect 114 31 116 33
rect 118 31 120 33
rect 114 29 120 31
rect 124 33 146 35
rect 124 31 135 33
rect 137 31 142 33
rect 144 31 146 33
rect 124 29 146 31
rect 150 33 156 35
rect 150 31 152 33
rect 154 31 156 33
rect 150 29 156 31
rect 160 33 166 35
rect 160 31 162 33
rect 164 31 166 33
rect 160 29 166 31
rect 182 33 188 35
rect 182 31 184 33
rect 186 31 188 33
rect 182 29 188 31
rect 192 33 198 35
rect 192 31 194 33
rect 196 31 198 33
rect 192 29 198 31
rect 202 33 224 35
rect 202 31 204 33
rect 206 31 211 33
rect 213 31 224 33
rect 202 29 224 31
rect 228 33 234 35
rect 228 31 230 33
rect 232 31 234 33
rect 228 29 234 31
rect 114 26 116 29
rect 124 26 126 29
rect 144 26 146 29
rect 151 26 153 29
rect 54 8 56 13
rect 61 8 63 13
rect 74 11 76 15
rect 94 2 96 6
rect 104 4 106 9
rect 114 7 116 12
rect 124 7 126 12
rect 162 20 164 29
rect 184 20 186 29
rect 195 26 197 29
rect 202 26 204 29
rect 222 26 224 29
rect 232 26 234 29
rect 242 34 244 36
rect 246 34 248 36
rect 242 32 248 34
rect 242 19 244 32
rect 252 28 254 41
rect 269 40 275 42
rect 269 38 271 40
rect 273 38 275 40
rect 269 36 275 38
rect 248 26 254 28
rect 273 26 275 36
rect 280 35 282 45
rect 341 57 343 61
rect 321 43 323 46
rect 317 41 323 43
rect 317 39 319 41
rect 321 39 323 41
rect 293 35 295 38
rect 317 37 323 39
rect 279 33 285 35
rect 279 31 281 33
rect 283 31 285 33
rect 279 29 285 31
rect 289 33 295 35
rect 289 31 291 33
rect 293 31 295 33
rect 289 29 295 31
rect 283 26 285 29
rect 293 26 295 29
rect 248 24 250 26
rect 252 24 254 26
rect 248 22 254 24
rect 252 19 254 22
rect 222 7 224 12
rect 232 7 234 12
rect 144 2 146 6
rect 151 2 153 6
rect 162 2 164 6
rect 184 2 186 6
rect 195 2 197 6
rect 202 2 204 6
rect 242 4 244 9
rect 273 15 275 20
rect 283 15 285 20
rect 321 24 323 37
rect 331 35 333 46
rect 394 63 396 68
rect 401 63 403 68
rect 419 66 421 70
rect 429 66 431 70
rect 439 66 441 70
rect 461 66 463 70
rect 471 66 473 70
rect 481 66 483 70
rect 384 54 386 59
rect 341 35 343 39
rect 327 33 333 35
rect 327 31 329 33
rect 331 31 333 33
rect 327 29 333 31
rect 337 33 343 35
rect 337 31 339 33
rect 341 31 343 33
rect 337 29 343 31
rect 328 24 330 29
rect 341 24 343 29
rect 371 28 373 41
rect 384 38 386 41
rect 499 63 501 68
rect 506 63 508 68
rect 529 66 531 70
rect 550 66 552 70
rect 557 66 559 70
rect 516 54 518 59
rect 647 66 649 70
rect 570 56 572 61
rect 598 59 600 64
rect 608 59 610 64
rect 550 42 552 45
rect 516 38 518 41
rect 377 36 386 38
rect 377 34 379 36
rect 381 34 383 36
rect 394 35 396 38
rect 401 35 403 38
rect 419 35 421 38
rect 429 35 431 38
rect 439 35 441 38
rect 461 35 463 38
rect 471 35 473 38
rect 481 35 483 38
rect 499 35 501 38
rect 506 35 508 38
rect 516 36 525 38
rect 377 32 383 34
rect 371 26 377 28
rect 371 24 373 26
rect 375 24 377 26
rect 293 12 295 17
rect 371 22 377 24
rect 371 19 373 22
rect 381 19 383 32
rect 391 33 397 35
rect 391 31 393 33
rect 395 31 397 33
rect 391 29 397 31
rect 401 33 423 35
rect 401 31 412 33
rect 414 31 419 33
rect 421 31 423 33
rect 401 29 423 31
rect 427 33 433 35
rect 427 31 429 33
rect 431 31 433 33
rect 427 29 433 31
rect 437 33 443 35
rect 437 31 439 33
rect 441 31 443 33
rect 437 29 443 31
rect 459 33 465 35
rect 459 31 461 33
rect 463 31 465 33
rect 459 29 465 31
rect 469 33 475 35
rect 469 31 471 33
rect 473 31 475 33
rect 469 29 475 31
rect 479 33 501 35
rect 479 31 481 33
rect 483 31 488 33
rect 490 31 501 33
rect 479 29 501 31
rect 505 33 511 35
rect 505 31 507 33
rect 509 31 511 33
rect 505 29 511 31
rect 391 26 393 29
rect 401 26 403 29
rect 421 26 423 29
rect 428 26 430 29
rect 321 8 323 13
rect 328 8 330 13
rect 252 2 254 6
rect 341 11 343 15
rect 371 2 373 6
rect 381 4 383 9
rect 391 7 393 12
rect 401 7 403 12
rect 439 20 441 29
rect 461 20 463 29
rect 472 26 474 29
rect 479 26 481 29
rect 499 26 501 29
rect 509 26 511 29
rect 519 34 521 36
rect 523 34 525 36
rect 519 32 525 34
rect 519 19 521 32
rect 529 28 531 41
rect 546 40 552 42
rect 546 38 548 40
rect 550 38 552 40
rect 546 36 552 38
rect 525 26 531 28
rect 550 26 552 36
rect 557 35 559 45
rect 618 57 620 61
rect 598 43 600 46
rect 594 41 600 43
rect 594 39 596 41
rect 598 39 600 41
rect 570 35 572 38
rect 594 37 600 39
rect 556 33 562 35
rect 556 31 558 33
rect 560 31 562 33
rect 556 29 562 31
rect 566 33 572 35
rect 566 31 568 33
rect 570 31 572 33
rect 566 29 572 31
rect 560 26 562 29
rect 570 26 572 29
rect 525 24 527 26
rect 529 24 531 26
rect 525 22 531 24
rect 529 19 531 22
rect 499 7 501 12
rect 509 7 511 12
rect 421 2 423 6
rect 428 2 430 6
rect 439 2 441 6
rect 461 2 463 6
rect 472 2 474 6
rect 479 2 481 6
rect 519 4 521 9
rect 550 15 552 20
rect 560 15 562 20
rect 598 24 600 37
rect 608 35 610 46
rect 670 63 672 68
rect 677 63 679 68
rect 695 66 697 70
rect 705 66 707 70
rect 715 66 717 70
rect 737 66 739 70
rect 747 66 749 70
rect 757 66 759 70
rect 660 54 662 59
rect 618 35 620 39
rect 604 33 610 35
rect 604 31 606 33
rect 608 31 610 33
rect 604 29 610 31
rect 614 33 620 35
rect 614 31 616 33
rect 618 31 620 33
rect 614 29 620 31
rect 605 24 607 29
rect 618 24 620 29
rect 647 28 649 41
rect 660 38 662 41
rect 775 63 777 68
rect 782 63 784 68
rect 805 66 807 70
rect 826 66 828 70
rect 833 66 835 70
rect 792 54 794 59
rect 924 66 926 70
rect 846 56 848 61
rect 874 59 876 64
rect 884 59 886 64
rect 826 42 828 45
rect 792 38 794 41
rect 653 36 662 38
rect 653 34 655 36
rect 657 34 659 36
rect 670 35 672 38
rect 677 35 679 38
rect 695 35 697 38
rect 705 35 707 38
rect 715 35 717 38
rect 737 35 739 38
rect 747 35 749 38
rect 757 35 759 38
rect 775 35 777 38
rect 782 35 784 38
rect 792 36 801 38
rect 653 32 659 34
rect 647 26 653 28
rect 647 24 649 26
rect 651 24 653 26
rect 570 12 572 17
rect 647 22 653 24
rect 647 19 649 22
rect 657 19 659 32
rect 667 33 673 35
rect 667 31 669 33
rect 671 31 673 33
rect 667 29 673 31
rect 677 33 699 35
rect 677 31 688 33
rect 690 31 695 33
rect 697 31 699 33
rect 677 29 699 31
rect 703 33 709 35
rect 703 31 705 33
rect 707 31 709 33
rect 703 29 709 31
rect 713 33 719 35
rect 713 31 715 33
rect 717 31 719 33
rect 713 29 719 31
rect 735 33 741 35
rect 735 31 737 33
rect 739 31 741 33
rect 735 29 741 31
rect 745 33 751 35
rect 745 31 747 33
rect 749 31 751 33
rect 745 29 751 31
rect 755 33 777 35
rect 755 31 757 33
rect 759 31 764 33
rect 766 31 777 33
rect 755 29 777 31
rect 781 33 787 35
rect 781 31 783 33
rect 785 31 787 33
rect 781 29 787 31
rect 667 26 669 29
rect 677 26 679 29
rect 697 26 699 29
rect 704 26 706 29
rect 598 8 600 13
rect 605 8 607 13
rect 529 2 531 6
rect 618 11 620 15
rect 647 2 649 6
rect 657 4 659 9
rect 667 7 669 12
rect 677 7 679 12
rect 715 20 717 29
rect 737 20 739 29
rect 748 26 750 29
rect 755 26 757 29
rect 775 26 777 29
rect 785 26 787 29
rect 795 34 797 36
rect 799 34 801 36
rect 795 32 801 34
rect 795 19 797 32
rect 805 28 807 41
rect 822 40 828 42
rect 822 38 824 40
rect 826 38 828 40
rect 822 36 828 38
rect 801 26 807 28
rect 826 26 828 36
rect 833 35 835 45
rect 894 57 896 61
rect 874 43 876 46
rect 870 41 876 43
rect 870 39 872 41
rect 874 39 876 41
rect 846 35 848 38
rect 870 37 876 39
rect 832 33 838 35
rect 832 31 834 33
rect 836 31 838 33
rect 832 29 838 31
rect 842 33 848 35
rect 842 31 844 33
rect 846 31 848 33
rect 842 29 848 31
rect 836 26 838 29
rect 846 26 848 29
rect 801 24 803 26
rect 805 24 807 26
rect 801 22 807 24
rect 805 19 807 22
rect 775 7 777 12
rect 785 7 787 12
rect 697 2 699 6
rect 704 2 706 6
rect 715 2 717 6
rect 737 2 739 6
rect 748 2 750 6
rect 755 2 757 6
rect 795 4 797 9
rect 826 15 828 20
rect 836 15 838 20
rect 874 24 876 37
rect 884 35 886 46
rect 947 63 949 68
rect 954 63 956 68
rect 972 66 974 70
rect 982 66 984 70
rect 992 66 994 70
rect 1014 66 1016 70
rect 1024 66 1026 70
rect 1034 66 1036 70
rect 937 54 939 59
rect 894 35 896 39
rect 880 33 886 35
rect 880 31 882 33
rect 884 31 886 33
rect 880 29 886 31
rect 890 33 896 35
rect 890 31 892 33
rect 894 31 896 33
rect 890 29 896 31
rect 881 24 883 29
rect 894 24 896 29
rect 924 28 926 41
rect 937 38 939 41
rect 1052 63 1054 68
rect 1059 63 1061 68
rect 1082 66 1084 70
rect 1103 66 1105 70
rect 1110 66 1112 70
rect 1069 54 1071 59
rect 1123 56 1125 61
rect 1103 42 1105 45
rect 1069 38 1071 41
rect 930 36 939 38
rect 930 34 932 36
rect 934 34 936 36
rect 947 35 949 38
rect 954 35 956 38
rect 972 35 974 38
rect 982 35 984 38
rect 992 35 994 38
rect 1014 35 1016 38
rect 1024 35 1026 38
rect 1034 35 1036 38
rect 1052 35 1054 38
rect 1059 35 1061 38
rect 1069 36 1078 38
rect 930 32 936 34
rect 924 26 930 28
rect 924 24 926 26
rect 928 24 930 26
rect 846 12 848 17
rect 924 22 930 24
rect 924 19 926 22
rect 934 19 936 32
rect 944 33 950 35
rect 944 31 946 33
rect 948 31 950 33
rect 944 29 950 31
rect 954 33 976 35
rect 954 31 965 33
rect 967 31 972 33
rect 974 31 976 33
rect 954 29 976 31
rect 980 33 986 35
rect 980 31 982 33
rect 984 31 986 33
rect 980 29 986 31
rect 990 33 996 35
rect 990 31 992 33
rect 994 31 996 33
rect 990 29 996 31
rect 1012 33 1018 35
rect 1012 31 1014 33
rect 1016 31 1018 33
rect 1012 29 1018 31
rect 1022 33 1028 35
rect 1022 31 1024 33
rect 1026 31 1028 33
rect 1022 29 1028 31
rect 1032 33 1054 35
rect 1032 31 1034 33
rect 1036 31 1041 33
rect 1043 31 1054 33
rect 1032 29 1054 31
rect 1058 33 1064 35
rect 1058 31 1060 33
rect 1062 31 1064 33
rect 1058 29 1064 31
rect 944 26 946 29
rect 954 26 956 29
rect 974 26 976 29
rect 981 26 983 29
rect 874 8 876 13
rect 881 8 883 13
rect 805 2 807 6
rect 894 11 896 15
rect 924 2 926 6
rect 934 4 936 9
rect 944 7 946 12
rect 954 7 956 12
rect 992 20 994 29
rect 1014 20 1016 29
rect 1025 26 1027 29
rect 1032 26 1034 29
rect 1052 26 1054 29
rect 1062 26 1064 29
rect 1072 34 1074 36
rect 1076 34 1078 36
rect 1072 32 1078 34
rect 1072 19 1074 32
rect 1082 28 1084 41
rect 1099 40 1105 42
rect 1099 38 1101 40
rect 1103 38 1105 40
rect 1099 36 1105 38
rect 1078 26 1084 28
rect 1103 26 1105 36
rect 1110 35 1112 45
rect 1123 35 1125 38
rect 1109 33 1115 35
rect 1109 31 1111 33
rect 1113 31 1115 33
rect 1109 29 1115 31
rect 1119 33 1125 35
rect 1119 31 1121 33
rect 1123 31 1125 33
rect 1119 29 1125 31
rect 1113 26 1115 29
rect 1123 26 1125 29
rect 1078 24 1080 26
rect 1082 24 1084 26
rect 1078 22 1084 24
rect 1082 19 1084 22
rect 1052 7 1054 12
rect 1062 7 1064 12
rect 974 2 976 6
rect 981 2 983 6
rect 992 2 994 6
rect 1014 2 1016 6
rect 1025 2 1027 6
rect 1032 2 1034 6
rect 1072 4 1074 9
rect 1103 15 1105 20
rect 1113 15 1115 20
rect 1123 12 1125 17
rect 1082 2 1084 6
rect -134 -14 -132 -9
rect -127 -14 -125 -9
rect -120 -14 -118 -10
rect -82 -14 -80 -9
rect -75 -14 -73 -9
rect -68 -14 -66 -10
rect -30 -14 -28 -9
rect -23 -14 -21 -9
rect -16 -14 -14 -10
rect 22 -14 24 -9
rect 29 -14 31 -9
rect 36 -14 38 -10
rect 74 -14 76 -9
rect 81 -14 83 -9
rect 88 -14 90 -10
rect 127 -14 129 -9
rect 134 -14 136 -9
rect 141 -14 143 -10
rect 315 -14 317 -9
rect 322 -14 324 -9
rect 329 -14 331 -10
rect 368 -14 370 -9
rect 375 -14 377 -9
rect 382 -14 384 -10
rect 420 -14 422 -9
rect 427 -14 429 -9
rect 434 -14 436 -10
rect 472 -14 474 -9
rect 479 -14 481 -9
rect 486 -14 488 -10
rect 524 -14 526 -9
rect 531 -14 533 -9
rect 538 -14 540 -10
rect 623 -14 625 -9
rect 630 -14 632 -9
rect 637 -14 639 -10
rect 676 -14 678 -9
rect 683 -14 685 -9
rect 690 -14 692 -10
rect 728 -14 730 -9
rect 735 -14 737 -9
rect 742 -14 744 -10
rect 780 -14 782 -9
rect 787 -14 789 -9
rect 794 -14 796 -10
rect 832 -14 834 -9
rect 839 -14 841 -9
rect 846 -14 848 -10
rect 884 -14 886 -9
rect 891 -14 893 -9
rect 898 -14 900 -10
rect 937 -14 939 -9
rect 944 -14 946 -9
rect 951 -14 953 -10
rect 991 -14 993 -9
rect 998 -14 1000 -9
rect 1005 -14 1007 -10
rect 1046 -14 1048 -9
rect 1053 -14 1055 -9
rect 1060 -14 1062 -10
rect 1099 -14 1101 -9
rect 1106 -14 1108 -9
rect 1113 -14 1115 -10
rect -149 -19 -147 -14
rect -97 -19 -95 -14
rect -45 -19 -43 -14
rect 7 -19 9 -14
rect 59 -19 61 -14
rect 112 -19 114 -14
rect 169 -19 171 -14
rect 189 -19 191 -14
rect 209 -19 211 -14
rect 231 -19 233 -14
rect 253 -19 255 -14
rect 275 -19 277 -14
rect 300 -19 302 -14
rect 353 -19 355 -14
rect 405 -19 407 -14
rect 457 -19 459 -14
rect 509 -19 511 -14
rect 564 -19 566 -14
rect 585 -19 587 -14
rect 608 -19 610 -14
rect 661 -19 663 -14
rect 713 -19 715 -14
rect 765 -19 767 -14
rect 817 -19 819 -14
rect 869 -19 871 -14
rect 922 -19 924 -14
rect 976 -19 978 -14
rect 1031 -19 1033 -14
rect 1084 -19 1086 -14
rect -149 -29 -147 -25
rect -134 -28 -132 -25
rect -149 -31 -143 -29
rect -149 -33 -147 -31
rect -145 -33 -143 -31
rect -149 -35 -143 -33
rect -139 -30 -132 -28
rect -139 -32 -137 -30
rect -135 -32 -132 -30
rect -139 -34 -132 -32
rect -149 -45 -147 -35
rect -139 -45 -137 -34
rect -127 -36 -125 -25
rect -120 -28 -118 -25
rect -120 -30 -111 -28
rect -117 -32 -115 -30
rect -113 -32 -111 -30
rect -117 -34 -111 -32
rect -97 -29 -95 -25
rect -82 -28 -80 -25
rect -97 -31 -91 -29
rect -97 -33 -95 -31
rect -93 -33 -91 -31
rect -127 -38 -121 -36
rect -127 -39 -125 -38
rect -129 -40 -125 -39
rect -123 -40 -121 -38
rect -129 -42 -121 -40
rect -129 -45 -127 -42
rect -117 -46 -115 -34
rect -97 -35 -91 -33
rect -87 -30 -80 -28
rect -87 -32 -85 -30
rect -83 -32 -80 -30
rect -87 -34 -80 -32
rect -97 -45 -95 -35
rect -87 -45 -85 -34
rect -75 -36 -73 -25
rect -68 -28 -66 -25
rect -68 -30 -59 -28
rect -65 -32 -63 -30
rect -61 -32 -59 -30
rect -65 -34 -59 -32
rect -45 -29 -43 -25
rect -30 -28 -28 -25
rect -45 -31 -39 -29
rect -45 -33 -43 -31
rect -41 -33 -39 -31
rect -75 -38 -69 -36
rect -75 -39 -73 -38
rect -77 -40 -73 -39
rect -71 -40 -69 -38
rect -77 -42 -69 -40
rect -77 -45 -75 -42
rect -149 -62 -147 -57
rect -139 -60 -137 -56
rect -129 -60 -127 -56
rect -65 -46 -63 -34
rect -45 -35 -39 -33
rect -35 -30 -28 -28
rect -35 -32 -33 -30
rect -31 -32 -28 -30
rect -35 -34 -28 -32
rect -45 -45 -43 -35
rect -35 -45 -33 -34
rect -23 -36 -21 -25
rect -16 -28 -14 -25
rect -16 -30 -7 -28
rect -13 -32 -11 -30
rect -9 -32 -7 -30
rect -13 -34 -7 -32
rect 7 -29 9 -25
rect 22 -28 24 -25
rect 7 -31 13 -29
rect 7 -33 9 -31
rect 11 -33 13 -31
rect -23 -38 -17 -36
rect -23 -39 -21 -38
rect -25 -40 -21 -39
rect -19 -40 -17 -38
rect -25 -42 -17 -40
rect -25 -45 -23 -42
rect -117 -61 -115 -57
rect -97 -62 -95 -57
rect -87 -60 -85 -56
rect -77 -60 -75 -56
rect -13 -46 -11 -34
rect 7 -35 13 -33
rect 17 -30 24 -28
rect 17 -32 19 -30
rect 21 -32 24 -30
rect 17 -34 24 -32
rect 7 -45 9 -35
rect 17 -45 19 -34
rect 29 -36 31 -25
rect 36 -28 38 -25
rect 36 -30 45 -28
rect 39 -32 41 -30
rect 43 -32 45 -30
rect 39 -34 45 -32
rect 59 -29 61 -25
rect 74 -28 76 -25
rect 59 -31 65 -29
rect 59 -33 61 -31
rect 63 -33 65 -31
rect 29 -38 35 -36
rect 29 -39 31 -38
rect 27 -40 31 -39
rect 33 -40 35 -38
rect 27 -42 35 -40
rect 27 -45 29 -42
rect -65 -61 -63 -57
rect -45 -62 -43 -57
rect -35 -60 -33 -56
rect -25 -60 -23 -56
rect 39 -46 41 -34
rect 59 -35 65 -33
rect 69 -30 76 -28
rect 69 -32 71 -30
rect 73 -32 76 -30
rect 69 -34 76 -32
rect 59 -45 61 -35
rect 69 -45 71 -34
rect 81 -36 83 -25
rect 88 -28 90 -25
rect 88 -30 97 -28
rect 91 -32 93 -30
rect 95 -32 97 -30
rect 91 -34 97 -32
rect 112 -29 114 -25
rect 127 -28 129 -25
rect 112 -31 118 -29
rect 112 -33 114 -31
rect 116 -33 118 -31
rect 81 -38 87 -36
rect 81 -39 83 -38
rect 79 -40 83 -39
rect 85 -40 87 -38
rect 79 -42 87 -40
rect 79 -45 81 -42
rect -13 -61 -11 -57
rect 7 -62 9 -57
rect 17 -60 19 -56
rect 27 -60 29 -56
rect 91 -46 93 -34
rect 112 -35 118 -33
rect 122 -30 129 -28
rect 122 -32 124 -30
rect 126 -32 129 -30
rect 122 -34 129 -32
rect 112 -45 114 -35
rect 122 -45 124 -34
rect 134 -36 136 -25
rect 141 -28 143 -25
rect 141 -30 150 -28
rect 144 -32 146 -30
rect 148 -32 150 -30
rect 144 -34 150 -32
rect 134 -38 140 -36
rect 134 -39 136 -38
rect 132 -40 136 -39
rect 138 -40 140 -38
rect 132 -42 140 -40
rect 132 -45 134 -42
rect 39 -61 41 -57
rect 59 -62 61 -57
rect 69 -60 71 -56
rect 79 -60 81 -56
rect 144 -46 146 -34
rect 169 -37 171 -25
rect 189 -37 191 -25
rect 209 -37 211 -25
rect 231 -37 233 -25
rect 253 -37 255 -25
rect 275 -37 277 -25
rect 300 -29 302 -25
rect 315 -28 317 -25
rect 300 -31 306 -29
rect 300 -33 302 -31
rect 304 -33 306 -31
rect 300 -35 306 -33
rect 310 -30 317 -28
rect 310 -32 312 -30
rect 314 -32 317 -30
rect 310 -34 317 -32
rect 91 -61 93 -57
rect 112 -62 114 -57
rect 122 -60 124 -56
rect 132 -60 134 -56
rect 300 -45 302 -35
rect 310 -45 312 -34
rect 322 -36 324 -25
rect 329 -28 331 -25
rect 329 -30 338 -28
rect 332 -32 334 -30
rect 336 -32 338 -30
rect 332 -34 338 -32
rect 353 -29 355 -25
rect 368 -28 370 -25
rect 353 -31 359 -29
rect 353 -33 355 -31
rect 357 -33 359 -31
rect 322 -38 328 -36
rect 322 -39 324 -38
rect 320 -40 324 -39
rect 326 -40 328 -38
rect 320 -42 328 -40
rect 320 -45 322 -42
rect 144 -61 146 -57
rect 169 -52 171 -49
rect 169 -54 175 -52
rect 169 -56 171 -54
rect 173 -56 175 -54
rect 169 -58 175 -56
rect 189 -52 191 -49
rect 189 -54 195 -52
rect 189 -56 191 -54
rect 193 -56 195 -54
rect 189 -58 195 -56
rect 209 -52 211 -49
rect 209 -54 215 -52
rect 209 -56 211 -54
rect 213 -56 215 -54
rect 209 -58 215 -56
rect 231 -52 233 -49
rect 231 -54 237 -52
rect 231 -56 233 -54
rect 235 -56 237 -54
rect 231 -58 237 -56
rect 253 -52 255 -49
rect 253 -54 259 -52
rect 253 -56 255 -54
rect 257 -56 259 -54
rect 253 -58 259 -56
rect 275 -52 277 -49
rect 275 -54 281 -52
rect 275 -56 277 -54
rect 279 -56 281 -54
rect 275 -58 281 -56
rect 332 -46 334 -34
rect 353 -35 359 -33
rect 363 -30 370 -28
rect 363 -32 365 -30
rect 367 -32 370 -30
rect 363 -34 370 -32
rect 353 -45 355 -35
rect 363 -45 365 -34
rect 375 -36 377 -25
rect 382 -28 384 -25
rect 382 -30 391 -28
rect 385 -32 387 -30
rect 389 -32 391 -30
rect 385 -34 391 -32
rect 405 -29 407 -25
rect 420 -28 422 -25
rect 405 -31 411 -29
rect 405 -33 407 -31
rect 409 -33 411 -31
rect 375 -38 381 -36
rect 375 -39 377 -38
rect 373 -40 377 -39
rect 379 -40 381 -38
rect 373 -42 381 -40
rect 373 -45 375 -42
rect 300 -62 302 -57
rect 310 -60 312 -56
rect 320 -60 322 -56
rect 385 -46 387 -34
rect 405 -35 411 -33
rect 415 -30 422 -28
rect 415 -32 417 -30
rect 419 -32 422 -30
rect 415 -34 422 -32
rect 405 -45 407 -35
rect 415 -45 417 -34
rect 427 -36 429 -25
rect 434 -28 436 -25
rect 434 -30 443 -28
rect 437 -32 439 -30
rect 441 -32 443 -30
rect 437 -34 443 -32
rect 457 -29 459 -25
rect 472 -28 474 -25
rect 457 -31 463 -29
rect 457 -33 459 -31
rect 461 -33 463 -31
rect 427 -38 433 -36
rect 427 -39 429 -38
rect 425 -40 429 -39
rect 431 -40 433 -38
rect 425 -42 433 -40
rect 425 -45 427 -42
rect 332 -61 334 -57
rect 353 -62 355 -57
rect 363 -60 365 -56
rect 373 -60 375 -56
rect 437 -46 439 -34
rect 457 -35 463 -33
rect 467 -30 474 -28
rect 467 -32 469 -30
rect 471 -32 474 -30
rect 467 -34 474 -32
rect 457 -45 459 -35
rect 467 -45 469 -34
rect 479 -36 481 -25
rect 486 -28 488 -25
rect 486 -30 495 -28
rect 489 -32 491 -30
rect 493 -32 495 -30
rect 489 -34 495 -32
rect 509 -29 511 -25
rect 524 -28 526 -25
rect 509 -31 515 -29
rect 509 -33 511 -31
rect 513 -33 515 -31
rect 479 -38 485 -36
rect 479 -39 481 -38
rect 477 -40 481 -39
rect 483 -40 485 -38
rect 477 -42 485 -40
rect 477 -45 479 -42
rect 385 -61 387 -57
rect 405 -62 407 -57
rect 415 -60 417 -56
rect 425 -60 427 -56
rect 489 -46 491 -34
rect 509 -35 515 -33
rect 519 -30 526 -28
rect 519 -32 521 -30
rect 523 -32 526 -30
rect 519 -34 526 -32
rect 509 -45 511 -35
rect 519 -45 521 -34
rect 531 -36 533 -25
rect 538 -28 540 -25
rect 538 -30 547 -28
rect 541 -32 543 -30
rect 545 -32 547 -30
rect 541 -34 547 -32
rect 531 -38 537 -36
rect 531 -39 533 -38
rect 529 -40 533 -39
rect 535 -40 537 -38
rect 529 -42 537 -40
rect 529 -45 531 -42
rect 437 -61 439 -57
rect 457 -62 459 -57
rect 467 -60 469 -56
rect 477 -60 479 -56
rect 541 -46 543 -34
rect 564 -37 566 -25
rect 585 -37 587 -25
rect 608 -29 610 -25
rect 623 -28 625 -25
rect 608 -31 614 -29
rect 608 -33 610 -31
rect 612 -33 614 -31
rect 608 -35 614 -33
rect 618 -30 625 -28
rect 618 -32 620 -30
rect 622 -32 625 -30
rect 618 -34 625 -32
rect 489 -61 491 -57
rect 509 -62 511 -57
rect 519 -60 521 -56
rect 529 -60 531 -56
rect 608 -45 610 -35
rect 618 -45 620 -34
rect 630 -36 632 -25
rect 637 -28 639 -25
rect 637 -30 646 -28
rect 640 -32 642 -30
rect 644 -32 646 -30
rect 640 -34 646 -32
rect 661 -29 663 -25
rect 676 -28 678 -25
rect 661 -31 667 -29
rect 661 -33 663 -31
rect 665 -33 667 -31
rect 630 -38 636 -36
rect 630 -39 632 -38
rect 628 -40 632 -39
rect 634 -40 636 -38
rect 628 -42 636 -40
rect 628 -45 630 -42
rect 541 -61 543 -57
rect 564 -52 566 -49
rect 564 -54 570 -52
rect 564 -56 566 -54
rect 568 -56 570 -54
rect 564 -58 570 -56
rect 585 -52 587 -49
rect 585 -54 591 -52
rect 585 -56 587 -54
rect 589 -56 591 -54
rect 585 -58 591 -56
rect 640 -46 642 -34
rect 661 -35 667 -33
rect 671 -30 678 -28
rect 671 -32 673 -30
rect 675 -32 678 -30
rect 671 -34 678 -32
rect 661 -45 663 -35
rect 671 -45 673 -34
rect 683 -36 685 -25
rect 690 -28 692 -25
rect 690 -30 699 -28
rect 693 -32 695 -30
rect 697 -32 699 -30
rect 693 -34 699 -32
rect 713 -29 715 -25
rect 728 -28 730 -25
rect 713 -31 719 -29
rect 713 -33 715 -31
rect 717 -33 719 -31
rect 683 -38 689 -36
rect 683 -39 685 -38
rect 681 -40 685 -39
rect 687 -40 689 -38
rect 681 -42 689 -40
rect 681 -45 683 -42
rect 608 -62 610 -57
rect 618 -60 620 -56
rect 628 -60 630 -56
rect 693 -46 695 -34
rect 713 -35 719 -33
rect 723 -30 730 -28
rect 723 -32 725 -30
rect 727 -32 730 -30
rect 723 -34 730 -32
rect 713 -45 715 -35
rect 723 -45 725 -34
rect 735 -36 737 -25
rect 742 -28 744 -25
rect 742 -30 751 -28
rect 745 -32 747 -30
rect 749 -32 751 -30
rect 745 -34 751 -32
rect 765 -29 767 -25
rect 780 -28 782 -25
rect 765 -31 771 -29
rect 765 -33 767 -31
rect 769 -33 771 -31
rect 735 -38 741 -36
rect 735 -39 737 -38
rect 733 -40 737 -39
rect 739 -40 741 -38
rect 733 -42 741 -40
rect 733 -45 735 -42
rect 640 -61 642 -57
rect 661 -62 663 -57
rect 671 -60 673 -56
rect 681 -60 683 -56
rect 745 -46 747 -34
rect 765 -35 771 -33
rect 775 -30 782 -28
rect 775 -32 777 -30
rect 779 -32 782 -30
rect 775 -34 782 -32
rect 765 -45 767 -35
rect 775 -45 777 -34
rect 787 -36 789 -25
rect 794 -28 796 -25
rect 794 -30 803 -28
rect 797 -32 799 -30
rect 801 -32 803 -30
rect 797 -34 803 -32
rect 817 -29 819 -25
rect 832 -28 834 -25
rect 817 -31 823 -29
rect 817 -33 819 -31
rect 821 -33 823 -31
rect 787 -38 793 -36
rect 787 -39 789 -38
rect 785 -40 789 -39
rect 791 -40 793 -38
rect 785 -42 793 -40
rect 785 -45 787 -42
rect 693 -61 695 -57
rect 713 -62 715 -57
rect 723 -60 725 -56
rect 733 -60 735 -56
rect 797 -46 799 -34
rect 817 -35 823 -33
rect 827 -30 834 -28
rect 827 -32 829 -30
rect 831 -32 834 -30
rect 827 -34 834 -32
rect 817 -45 819 -35
rect 827 -45 829 -34
rect 839 -36 841 -25
rect 846 -28 848 -25
rect 846 -30 855 -28
rect 849 -32 851 -30
rect 853 -32 855 -30
rect 849 -34 855 -32
rect 869 -29 871 -25
rect 884 -28 886 -25
rect 869 -31 875 -29
rect 869 -33 871 -31
rect 873 -33 875 -31
rect 839 -38 845 -36
rect 839 -39 841 -38
rect 837 -40 841 -39
rect 843 -40 845 -38
rect 837 -42 845 -40
rect 837 -45 839 -42
rect 745 -61 747 -57
rect 765 -62 767 -57
rect 775 -60 777 -56
rect 785 -60 787 -56
rect 849 -46 851 -34
rect 869 -35 875 -33
rect 879 -30 886 -28
rect 879 -32 881 -30
rect 883 -32 886 -30
rect 879 -34 886 -32
rect 869 -45 871 -35
rect 879 -45 881 -34
rect 891 -36 893 -25
rect 898 -28 900 -25
rect 898 -30 907 -28
rect 901 -32 903 -30
rect 905 -32 907 -30
rect 901 -34 907 -32
rect 922 -29 924 -25
rect 937 -28 939 -25
rect 922 -31 928 -29
rect 922 -33 924 -31
rect 926 -33 928 -31
rect 891 -38 897 -36
rect 891 -39 893 -38
rect 889 -40 893 -39
rect 895 -40 897 -38
rect 889 -42 897 -40
rect 889 -45 891 -42
rect 797 -61 799 -57
rect 817 -62 819 -57
rect 827 -60 829 -56
rect 837 -60 839 -56
rect 901 -46 903 -34
rect 922 -35 928 -33
rect 932 -30 939 -28
rect 932 -32 934 -30
rect 936 -32 939 -30
rect 932 -34 939 -32
rect 922 -45 924 -35
rect 932 -45 934 -34
rect 944 -36 946 -25
rect 951 -28 953 -25
rect 951 -30 960 -28
rect 954 -32 956 -30
rect 958 -32 960 -30
rect 954 -34 960 -32
rect 976 -29 978 -25
rect 991 -28 993 -25
rect 976 -31 982 -29
rect 976 -33 978 -31
rect 980 -33 982 -31
rect 944 -38 950 -36
rect 944 -39 946 -38
rect 942 -40 946 -39
rect 948 -40 950 -38
rect 942 -42 950 -40
rect 942 -45 944 -42
rect 849 -61 851 -57
rect 869 -62 871 -57
rect 879 -60 881 -56
rect 889 -60 891 -56
rect 954 -46 956 -34
rect 976 -35 982 -33
rect 986 -30 993 -28
rect 986 -32 988 -30
rect 990 -32 993 -30
rect 986 -34 993 -32
rect 976 -45 978 -35
rect 986 -45 988 -34
rect 998 -36 1000 -25
rect 1005 -28 1007 -25
rect 1005 -30 1014 -28
rect 1008 -32 1010 -30
rect 1012 -32 1014 -30
rect 1008 -34 1014 -32
rect 1031 -29 1033 -25
rect 1046 -28 1048 -25
rect 1031 -31 1037 -29
rect 1031 -33 1033 -31
rect 1035 -33 1037 -31
rect 998 -38 1004 -36
rect 998 -39 1000 -38
rect 996 -40 1000 -39
rect 1002 -40 1004 -38
rect 996 -42 1004 -40
rect 996 -45 998 -42
rect 901 -61 903 -57
rect 922 -62 924 -57
rect 932 -60 934 -56
rect 942 -60 944 -56
rect 1008 -46 1010 -34
rect 1031 -35 1037 -33
rect 1041 -30 1048 -28
rect 1041 -32 1043 -30
rect 1045 -32 1048 -30
rect 1041 -34 1048 -32
rect 1031 -45 1033 -35
rect 1041 -45 1043 -34
rect 1053 -36 1055 -25
rect 1060 -28 1062 -25
rect 1060 -30 1069 -28
rect 1063 -32 1065 -30
rect 1067 -32 1069 -30
rect 1063 -34 1069 -32
rect 1084 -29 1086 -25
rect 1099 -28 1101 -25
rect 1084 -31 1090 -29
rect 1084 -33 1086 -31
rect 1088 -33 1090 -31
rect 1053 -38 1059 -36
rect 1053 -39 1055 -38
rect 1051 -40 1055 -39
rect 1057 -40 1059 -38
rect 1051 -42 1059 -40
rect 1051 -45 1053 -42
rect 954 -61 956 -57
rect 976 -62 978 -57
rect 986 -60 988 -56
rect 996 -60 998 -56
rect 1063 -46 1065 -34
rect 1084 -35 1090 -33
rect 1094 -30 1101 -28
rect 1094 -32 1096 -30
rect 1098 -32 1101 -30
rect 1094 -34 1101 -32
rect 1084 -45 1086 -35
rect 1094 -45 1096 -34
rect 1106 -36 1108 -25
rect 1113 -28 1115 -25
rect 1113 -30 1122 -28
rect 1116 -32 1118 -30
rect 1120 -32 1122 -30
rect 1116 -34 1122 -32
rect 1106 -38 1112 -36
rect 1106 -39 1108 -38
rect 1104 -40 1108 -39
rect 1110 -40 1112 -38
rect 1104 -42 1112 -40
rect 1104 -45 1106 -42
rect 1008 -61 1010 -57
rect 1031 -62 1033 -57
rect 1041 -60 1043 -56
rect 1051 -60 1053 -56
rect 1116 -46 1118 -34
rect 1063 -61 1065 -57
rect 1084 -62 1086 -57
rect 1094 -60 1096 -56
rect 1104 -60 1106 -56
rect 1116 -61 1118 -57
<< ndif >>
rect -283 312 -276 314
rect -283 310 -281 312
rect -279 310 -276 312
rect -283 308 -276 310
rect -281 305 -276 308
rect -274 309 -269 314
rect -274 305 -260 309
rect -269 304 -260 305
rect -269 302 -267 304
rect -265 302 -260 304
rect -269 300 -260 302
rect -258 307 -250 309
rect -258 305 -255 307
rect -253 305 -250 307
rect -258 300 -250 305
rect -248 305 -240 309
rect -248 303 -245 305
rect -243 303 -240 305
rect -248 300 -240 303
rect -245 297 -240 300
rect -238 297 -233 309
rect -231 297 -223 309
rect -193 307 -188 314
rect -215 305 -208 307
rect -215 303 -213 305
rect -211 303 -208 305
rect -215 301 -208 303
rect -229 295 -223 297
rect -229 293 -227 295
rect -225 293 -223 295
rect -213 294 -208 301
rect -206 301 -198 307
rect -206 299 -203 301
rect -201 299 -198 301
rect -206 297 -198 299
rect -196 304 -188 307
rect -196 302 -193 304
rect -191 302 -188 304
rect -196 300 -188 302
rect -186 312 -178 314
rect -186 310 -183 312
rect -181 310 -178 312
rect -186 300 -178 310
rect -176 312 -169 314
rect -176 310 -173 312
rect -171 310 -169 312
rect -176 305 -169 310
rect -163 307 -158 314
rect -176 303 -173 305
rect -171 303 -169 305
rect -176 300 -169 303
rect -165 305 -158 307
rect -165 303 -163 305
rect -161 303 -158 305
rect -165 301 -158 303
rect -196 297 -191 300
rect -206 294 -201 297
rect -229 291 -223 293
rect -163 294 -158 301
rect -156 294 -151 314
rect -149 308 -142 314
rect -114 308 -107 314
rect -149 298 -140 308
rect -149 296 -146 298
rect -144 296 -140 298
rect -149 294 -140 296
rect -138 305 -131 308
rect -138 303 -135 305
rect -133 303 -131 305
rect -138 301 -131 303
rect -125 305 -118 308
rect -125 303 -123 305
rect -121 303 -118 305
rect -125 301 -118 303
rect -138 294 -133 301
rect -123 294 -118 301
rect -116 298 -107 308
rect -116 296 -112 298
rect -110 296 -107 298
rect -116 294 -107 296
rect -105 294 -100 314
rect -98 307 -93 314
rect -87 312 -80 314
rect -87 310 -85 312
rect -83 310 -80 312
rect -98 305 -91 307
rect -98 303 -95 305
rect -93 303 -91 305
rect -98 301 -91 303
rect -87 305 -80 310
rect -87 303 -85 305
rect -83 303 -80 305
rect -98 294 -93 301
rect -87 300 -80 303
rect -78 312 -70 314
rect -78 310 -75 312
rect -73 310 -70 312
rect -78 300 -70 310
rect -68 307 -63 314
rect -36 308 -29 314
rect -27 312 -19 314
rect -27 310 -24 312
rect -22 310 -19 312
rect -27 308 -19 310
rect -17 308 -9 314
rect -68 304 -60 307
rect -68 302 -65 304
rect -63 302 -60 304
rect -68 300 -60 302
rect -65 297 -60 300
rect -58 301 -50 307
rect -58 299 -55 301
rect -53 299 -50 301
rect -58 297 -50 299
rect -55 294 -50 297
rect -48 305 -41 307
rect -48 303 -45 305
rect -43 303 -41 305
rect -48 301 -41 303
rect -36 301 -31 308
rect -15 305 -9 308
rect -7 312 0 314
rect -7 310 -4 312
rect -2 310 0 312
rect -7 308 0 310
rect -7 305 -2 308
rect 9 307 14 312
rect 7 305 14 307
rect -15 301 -11 305
rect -48 294 -43 301
rect -36 299 -30 301
rect -36 297 -34 299
rect -32 297 -30 299
rect -36 295 -30 297
rect -17 299 -11 301
rect 7 303 9 305
rect 11 303 14 305
rect 7 301 14 303
rect 16 301 21 312
rect 23 303 34 312
rect 36 309 41 312
rect 36 307 43 309
rect 49 307 54 312
rect 36 305 39 307
rect 41 305 43 307
rect 36 303 43 305
rect 47 305 54 307
rect 47 303 49 305
rect 51 303 54 305
rect 23 301 32 303
rect -17 297 -15 299
rect -13 297 -11 299
rect -17 295 -11 297
rect 25 295 32 301
rect 47 301 54 303
rect 56 301 61 312
rect 63 303 74 312
rect 76 309 81 312
rect 76 307 83 309
rect 109 307 114 314
rect 76 305 79 307
rect 81 305 83 307
rect 76 303 83 305
rect 87 305 94 307
rect 87 303 89 305
rect 91 303 94 305
rect 63 301 72 303
rect 25 293 28 295
rect 30 293 32 295
rect 25 291 32 293
rect 65 295 72 301
rect 87 301 94 303
rect 65 293 68 295
rect 70 293 72 295
rect 65 291 72 293
rect 89 294 94 301
rect 96 301 104 307
rect 96 299 99 301
rect 101 299 104 301
rect 96 297 104 299
rect 106 304 114 307
rect 106 302 109 304
rect 111 302 114 304
rect 106 300 114 302
rect 116 312 124 314
rect 116 310 119 312
rect 121 310 124 312
rect 116 300 124 310
rect 126 312 133 314
rect 126 310 129 312
rect 131 310 133 312
rect 126 305 133 310
rect 139 307 144 314
rect 126 303 129 305
rect 131 303 133 305
rect 126 300 133 303
rect 137 305 144 307
rect 137 303 139 305
rect 141 303 144 305
rect 137 301 144 303
rect 106 297 111 300
rect 96 294 101 297
rect 139 294 144 301
rect 146 294 151 314
rect 153 308 160 314
rect 188 308 195 314
rect 153 298 162 308
rect 153 296 156 298
rect 158 296 162 298
rect 153 294 162 296
rect 164 305 171 308
rect 164 303 167 305
rect 169 303 171 305
rect 164 301 171 303
rect 177 305 184 308
rect 177 303 179 305
rect 181 303 184 305
rect 177 301 184 303
rect 164 294 169 301
rect 179 294 184 301
rect 186 298 195 308
rect 186 296 190 298
rect 192 296 195 298
rect 186 294 195 296
rect 197 294 202 314
rect 204 307 209 314
rect 215 312 222 314
rect 215 310 217 312
rect 219 310 222 312
rect 204 305 211 307
rect 204 303 207 305
rect 209 303 211 305
rect 204 301 211 303
rect 215 305 222 310
rect 215 303 217 305
rect 219 303 222 305
rect 204 294 209 301
rect 215 300 222 303
rect 224 312 232 314
rect 224 310 227 312
rect 229 310 232 312
rect 224 300 232 310
rect 234 307 239 314
rect 266 308 273 314
rect 275 312 283 314
rect 275 310 278 312
rect 280 310 283 312
rect 275 308 283 310
rect 285 308 293 314
rect 234 304 242 307
rect 234 302 237 304
rect 239 302 242 304
rect 234 300 242 302
rect 237 297 242 300
rect 244 301 252 307
rect 244 299 247 301
rect 249 299 252 301
rect 244 297 252 299
rect 247 294 252 297
rect 254 305 261 307
rect 254 303 257 305
rect 259 303 261 305
rect 254 301 261 303
rect 266 301 271 308
rect 287 305 293 308
rect 295 312 302 314
rect 295 310 298 312
rect 300 310 302 312
rect 295 308 302 310
rect 295 305 300 308
rect 316 307 321 312
rect 314 305 321 307
rect 287 301 291 305
rect 254 294 259 301
rect 266 299 272 301
rect 266 297 268 299
rect 270 297 272 299
rect 266 295 272 297
rect 285 299 291 301
rect 314 303 316 305
rect 318 303 321 305
rect 314 301 321 303
rect 323 301 328 312
rect 330 303 341 312
rect 343 309 348 312
rect 343 307 350 309
rect 386 307 391 314
rect 343 305 346 307
rect 348 305 350 307
rect 343 303 350 305
rect 364 305 371 307
rect 364 303 366 305
rect 368 303 371 305
rect 330 301 339 303
rect 285 297 287 299
rect 289 297 291 299
rect 285 295 291 297
rect 332 295 339 301
rect 364 301 371 303
rect 332 293 335 295
rect 337 293 339 295
rect 332 291 339 293
rect 366 294 371 301
rect 373 301 381 307
rect 373 299 376 301
rect 378 299 381 301
rect 373 297 381 299
rect 383 304 391 307
rect 383 302 386 304
rect 388 302 391 304
rect 383 300 391 302
rect 393 312 401 314
rect 393 310 396 312
rect 398 310 401 312
rect 393 300 401 310
rect 403 312 410 314
rect 403 310 406 312
rect 408 310 410 312
rect 403 305 410 310
rect 416 307 421 314
rect 403 303 406 305
rect 408 303 410 305
rect 403 300 410 303
rect 414 305 421 307
rect 414 303 416 305
rect 418 303 421 305
rect 414 301 421 303
rect 383 297 388 300
rect 373 294 378 297
rect 416 294 421 301
rect 423 294 428 314
rect 430 308 437 314
rect 465 308 472 314
rect 430 298 439 308
rect 430 296 433 298
rect 435 296 439 298
rect 430 294 439 296
rect 441 305 448 308
rect 441 303 444 305
rect 446 303 448 305
rect 441 301 448 303
rect 454 305 461 308
rect 454 303 456 305
rect 458 303 461 305
rect 454 301 461 303
rect 441 294 446 301
rect 456 294 461 301
rect 463 298 472 308
rect 463 296 467 298
rect 469 296 472 298
rect 463 294 472 296
rect 474 294 479 314
rect 481 307 486 314
rect 492 312 499 314
rect 492 310 494 312
rect 496 310 499 312
rect 481 305 488 307
rect 481 303 484 305
rect 486 303 488 305
rect 481 301 488 303
rect 492 305 499 310
rect 492 303 494 305
rect 496 303 499 305
rect 481 294 486 301
rect 492 300 499 303
rect 501 312 509 314
rect 501 310 504 312
rect 506 310 509 312
rect 501 300 509 310
rect 511 307 516 314
rect 543 308 550 314
rect 552 312 560 314
rect 552 310 555 312
rect 557 310 560 312
rect 552 308 560 310
rect 562 308 570 314
rect 511 304 519 307
rect 511 302 514 304
rect 516 302 519 304
rect 511 300 519 302
rect 514 297 519 300
rect 521 301 529 307
rect 521 299 524 301
rect 526 299 529 301
rect 521 297 529 299
rect 524 294 529 297
rect 531 305 538 307
rect 531 303 534 305
rect 536 303 538 305
rect 531 301 538 303
rect 543 301 548 308
rect 564 305 570 308
rect 572 312 579 314
rect 572 310 575 312
rect 577 310 579 312
rect 572 308 579 310
rect 572 305 577 308
rect 593 307 598 312
rect 591 305 598 307
rect 564 301 568 305
rect 531 294 536 301
rect 543 299 549 301
rect 543 297 545 299
rect 547 297 549 299
rect 543 295 549 297
rect 562 299 568 301
rect 591 303 593 305
rect 595 303 598 305
rect 591 301 598 303
rect 600 301 605 312
rect 607 303 618 312
rect 620 309 625 312
rect 620 307 627 309
rect 662 307 667 314
rect 620 305 623 307
rect 625 305 627 307
rect 620 303 627 305
rect 640 305 647 307
rect 640 303 642 305
rect 644 303 647 305
rect 607 301 616 303
rect 562 297 564 299
rect 566 297 568 299
rect 562 295 568 297
rect 609 295 616 301
rect 640 301 647 303
rect 609 293 612 295
rect 614 293 616 295
rect 609 291 616 293
rect 642 294 647 301
rect 649 301 657 307
rect 649 299 652 301
rect 654 299 657 301
rect 649 297 657 299
rect 659 304 667 307
rect 659 302 662 304
rect 664 302 667 304
rect 659 300 667 302
rect 669 312 677 314
rect 669 310 672 312
rect 674 310 677 312
rect 669 300 677 310
rect 679 312 686 314
rect 679 310 682 312
rect 684 310 686 312
rect 679 305 686 310
rect 692 307 697 314
rect 679 303 682 305
rect 684 303 686 305
rect 679 300 686 303
rect 690 305 697 307
rect 690 303 692 305
rect 694 303 697 305
rect 690 301 697 303
rect 659 297 664 300
rect 649 294 654 297
rect 692 294 697 301
rect 699 294 704 314
rect 706 308 713 314
rect 741 308 748 314
rect 706 298 715 308
rect 706 296 709 298
rect 711 296 715 298
rect 706 294 715 296
rect 717 305 724 308
rect 717 303 720 305
rect 722 303 724 305
rect 717 301 724 303
rect 730 305 737 308
rect 730 303 732 305
rect 734 303 737 305
rect 730 301 737 303
rect 717 294 722 301
rect 732 294 737 301
rect 739 298 748 308
rect 739 296 743 298
rect 745 296 748 298
rect 739 294 748 296
rect 750 294 755 314
rect 757 307 762 314
rect 768 312 775 314
rect 768 310 770 312
rect 772 310 775 312
rect 757 305 764 307
rect 757 303 760 305
rect 762 303 764 305
rect 757 301 764 303
rect 768 305 775 310
rect 768 303 770 305
rect 772 303 775 305
rect 757 294 762 301
rect 768 300 775 303
rect 777 312 785 314
rect 777 310 780 312
rect 782 310 785 312
rect 777 300 785 310
rect 787 307 792 314
rect 819 308 826 314
rect 828 312 836 314
rect 828 310 831 312
rect 833 310 836 312
rect 828 308 836 310
rect 838 308 846 314
rect 787 304 795 307
rect 787 302 790 304
rect 792 302 795 304
rect 787 300 795 302
rect 790 297 795 300
rect 797 301 805 307
rect 797 299 800 301
rect 802 299 805 301
rect 797 297 805 299
rect 800 294 805 297
rect 807 305 814 307
rect 807 303 810 305
rect 812 303 814 305
rect 807 301 814 303
rect 819 301 824 308
rect 840 305 846 308
rect 848 312 855 314
rect 848 310 851 312
rect 853 310 855 312
rect 848 308 855 310
rect 848 305 853 308
rect 869 307 874 312
rect 867 305 874 307
rect 840 301 844 305
rect 807 294 812 301
rect 819 299 825 301
rect 819 297 821 299
rect 823 297 825 299
rect 819 295 825 297
rect 838 299 844 301
rect 867 303 869 305
rect 871 303 874 305
rect 867 301 874 303
rect 876 301 881 312
rect 883 303 894 312
rect 896 309 901 312
rect 896 307 903 309
rect 939 307 944 314
rect 896 305 899 307
rect 901 305 903 307
rect 896 303 903 305
rect 917 305 924 307
rect 917 303 919 305
rect 921 303 924 305
rect 883 301 892 303
rect 838 297 840 299
rect 842 297 844 299
rect 838 295 844 297
rect 885 295 892 301
rect 917 301 924 303
rect 885 293 888 295
rect 890 293 892 295
rect 885 291 892 293
rect 919 294 924 301
rect 926 301 934 307
rect 926 299 929 301
rect 931 299 934 301
rect 926 297 934 299
rect 936 304 944 307
rect 936 302 939 304
rect 941 302 944 304
rect 936 300 944 302
rect 946 312 954 314
rect 946 310 949 312
rect 951 310 954 312
rect 946 300 954 310
rect 956 312 963 314
rect 956 310 959 312
rect 961 310 963 312
rect 956 305 963 310
rect 969 307 974 314
rect 956 303 959 305
rect 961 303 963 305
rect 956 300 963 303
rect 967 305 974 307
rect 967 303 969 305
rect 971 303 974 305
rect 967 301 974 303
rect 936 297 941 300
rect 926 294 931 297
rect 969 294 974 301
rect 976 294 981 314
rect 983 308 990 314
rect 1018 308 1025 314
rect 983 298 992 308
rect 983 296 986 298
rect 988 296 992 298
rect 983 294 992 296
rect 994 305 1001 308
rect 994 303 997 305
rect 999 303 1001 305
rect 994 301 1001 303
rect 1007 305 1014 308
rect 1007 303 1009 305
rect 1011 303 1014 305
rect 1007 301 1014 303
rect 994 294 999 301
rect 1009 294 1014 301
rect 1016 298 1025 308
rect 1016 296 1020 298
rect 1022 296 1025 298
rect 1016 294 1025 296
rect 1027 294 1032 314
rect 1034 307 1039 314
rect 1045 312 1052 314
rect 1045 310 1047 312
rect 1049 310 1052 312
rect 1034 305 1041 307
rect 1034 303 1037 305
rect 1039 303 1041 305
rect 1034 301 1041 303
rect 1045 305 1052 310
rect 1045 303 1047 305
rect 1049 303 1052 305
rect 1034 294 1039 301
rect 1045 300 1052 303
rect 1054 312 1062 314
rect 1054 310 1057 312
rect 1059 310 1062 312
rect 1054 300 1062 310
rect 1064 307 1069 314
rect 1096 308 1103 314
rect 1105 312 1113 314
rect 1105 310 1108 312
rect 1110 310 1113 312
rect 1105 308 1113 310
rect 1115 308 1123 314
rect 1064 304 1072 307
rect 1064 302 1067 304
rect 1069 302 1072 304
rect 1064 300 1072 302
rect 1067 297 1072 300
rect 1074 301 1082 307
rect 1074 299 1077 301
rect 1079 299 1082 301
rect 1074 297 1082 299
rect 1077 294 1082 297
rect 1084 305 1091 307
rect 1084 303 1087 305
rect 1089 303 1091 305
rect 1084 301 1091 303
rect 1096 301 1101 308
rect 1117 305 1123 308
rect 1125 312 1132 314
rect 1125 310 1128 312
rect 1130 310 1132 312
rect 1125 308 1132 310
rect 1125 305 1130 308
rect 1117 301 1121 305
rect 1084 294 1089 301
rect 1096 299 1102 301
rect 1096 297 1098 299
rect 1100 297 1102 299
rect 1096 295 1102 297
rect 1115 299 1121 301
rect 1115 297 1117 299
rect 1119 297 1121 299
rect 1115 295 1121 297
rect -229 283 -223 285
rect -229 281 -227 283
rect -225 281 -223 283
rect -229 279 -223 281
rect -245 276 -240 279
rect -269 274 -260 276
rect -269 272 -267 274
rect -265 272 -260 274
rect -269 271 -260 272
rect -281 268 -276 271
rect -283 266 -276 268
rect -283 264 -281 266
rect -279 264 -276 266
rect -283 262 -276 264
rect -274 267 -260 271
rect -258 271 -250 276
rect -258 269 -255 271
rect -253 269 -250 271
rect -258 267 -250 269
rect -248 273 -240 276
rect -248 271 -245 273
rect -243 271 -240 273
rect -248 267 -240 271
rect -238 267 -233 279
rect -231 267 -223 279
rect -213 275 -208 282
rect -215 273 -208 275
rect -215 271 -213 273
rect -211 271 -208 273
rect -215 269 -208 271
rect -206 279 -201 282
rect -206 277 -198 279
rect -206 275 -203 277
rect -201 275 -198 277
rect -206 269 -198 275
rect -196 276 -191 279
rect -196 274 -188 276
rect -196 272 -193 274
rect -191 272 -188 274
rect -196 269 -188 272
rect -274 262 -269 267
rect -193 262 -188 269
rect -186 266 -178 276
rect -186 264 -183 266
rect -181 264 -178 266
rect -186 262 -178 264
rect -176 273 -169 276
rect -163 275 -158 282
rect -176 271 -173 273
rect -171 271 -169 273
rect -176 266 -169 271
rect -165 273 -158 275
rect -165 271 -163 273
rect -161 271 -158 273
rect -165 269 -158 271
rect -176 264 -173 266
rect -171 264 -169 266
rect -176 262 -169 264
rect -163 262 -158 269
rect -156 262 -151 282
rect -149 280 -140 282
rect -149 278 -146 280
rect -144 278 -140 280
rect -149 268 -140 278
rect -138 275 -133 282
rect -123 275 -118 282
rect -138 273 -131 275
rect -138 271 -135 273
rect -133 271 -131 273
rect -138 268 -131 271
rect -125 273 -118 275
rect -125 271 -123 273
rect -121 271 -118 273
rect -125 268 -118 271
rect -116 280 -107 282
rect -116 278 -112 280
rect -110 278 -107 280
rect -116 268 -107 278
rect -149 262 -142 268
rect -114 262 -107 268
rect -105 262 -100 282
rect -98 275 -93 282
rect -55 279 -50 282
rect -65 276 -60 279
rect -98 273 -91 275
rect -98 271 -95 273
rect -93 271 -91 273
rect -98 269 -91 271
rect -87 273 -80 276
rect -87 271 -85 273
rect -83 271 -80 273
rect -98 262 -93 269
rect -87 266 -80 271
rect -87 264 -85 266
rect -83 264 -80 266
rect -87 262 -80 264
rect -78 266 -70 276
rect -78 264 -75 266
rect -73 264 -70 266
rect -78 262 -70 264
rect -68 274 -60 276
rect -68 272 -65 274
rect -63 272 -60 274
rect -68 269 -60 272
rect -58 277 -50 279
rect -58 275 -55 277
rect -53 275 -50 277
rect -58 269 -50 275
rect -48 275 -43 282
rect -36 279 -30 281
rect -36 277 -34 279
rect -32 277 -30 279
rect -36 275 -30 277
rect -17 279 -11 281
rect 25 283 32 285
rect 25 281 28 283
rect 30 281 32 283
rect -17 277 -15 279
rect -13 277 -11 279
rect -17 275 -11 277
rect -48 273 -41 275
rect -48 271 -45 273
rect -43 271 -41 273
rect -48 269 -41 271
rect -68 262 -63 269
rect -36 268 -31 275
rect -15 271 -11 275
rect 25 275 32 281
rect 65 283 72 285
rect 65 281 68 283
rect 70 281 72 283
rect 7 273 14 275
rect 7 271 9 273
rect 11 271 14 273
rect -15 268 -9 271
rect -36 262 -29 268
rect -27 266 -19 268
rect -27 264 -24 266
rect -22 264 -19 266
rect -27 262 -19 264
rect -17 262 -9 268
rect -7 268 -2 271
rect 7 269 14 271
rect -7 266 0 268
rect -7 264 -4 266
rect -2 264 0 266
rect 9 264 14 269
rect 16 264 21 275
rect 23 273 32 275
rect 65 275 72 281
rect 47 273 54 275
rect 23 264 34 273
rect 36 271 43 273
rect 36 269 39 271
rect 41 269 43 271
rect 47 271 49 273
rect 51 271 54 273
rect 47 269 54 271
rect 36 267 43 269
rect 36 264 41 267
rect 49 264 54 269
rect 56 264 61 275
rect 63 273 72 275
rect 89 275 94 282
rect 87 273 94 275
rect 63 264 74 273
rect 76 271 83 273
rect 76 269 79 271
rect 81 269 83 271
rect 87 271 89 273
rect 91 271 94 273
rect 87 269 94 271
rect 96 279 101 282
rect 96 277 104 279
rect 96 275 99 277
rect 101 275 104 277
rect 96 269 104 275
rect 106 276 111 279
rect 106 274 114 276
rect 106 272 109 274
rect 111 272 114 274
rect 106 269 114 272
rect 76 267 83 269
rect 76 264 81 267
rect -7 262 0 264
rect 109 262 114 269
rect 116 266 124 276
rect 116 264 119 266
rect 121 264 124 266
rect 116 262 124 264
rect 126 273 133 276
rect 139 275 144 282
rect 126 271 129 273
rect 131 271 133 273
rect 126 266 133 271
rect 137 273 144 275
rect 137 271 139 273
rect 141 271 144 273
rect 137 269 144 271
rect 126 264 129 266
rect 131 264 133 266
rect 126 262 133 264
rect 139 262 144 269
rect 146 262 151 282
rect 153 280 162 282
rect 153 278 156 280
rect 158 278 162 280
rect 153 268 162 278
rect 164 275 169 282
rect 179 275 184 282
rect 164 273 171 275
rect 164 271 167 273
rect 169 271 171 273
rect 164 268 171 271
rect 177 273 184 275
rect 177 271 179 273
rect 181 271 184 273
rect 177 268 184 271
rect 186 280 195 282
rect 186 278 190 280
rect 192 278 195 280
rect 186 268 195 278
rect 153 262 160 268
rect 188 262 195 268
rect 197 262 202 282
rect 204 275 209 282
rect 247 279 252 282
rect 237 276 242 279
rect 204 273 211 275
rect 204 271 207 273
rect 209 271 211 273
rect 204 269 211 271
rect 215 273 222 276
rect 215 271 217 273
rect 219 271 222 273
rect 204 262 209 269
rect 215 266 222 271
rect 215 264 217 266
rect 219 264 222 266
rect 215 262 222 264
rect 224 266 232 276
rect 224 264 227 266
rect 229 264 232 266
rect 224 262 232 264
rect 234 274 242 276
rect 234 272 237 274
rect 239 272 242 274
rect 234 269 242 272
rect 244 277 252 279
rect 244 275 247 277
rect 249 275 252 277
rect 244 269 252 275
rect 254 275 259 282
rect 266 279 272 281
rect 266 277 268 279
rect 270 277 272 279
rect 266 275 272 277
rect 285 279 291 281
rect 332 283 339 285
rect 332 281 335 283
rect 337 281 339 283
rect 285 277 287 279
rect 289 277 291 279
rect 285 275 291 277
rect 254 273 261 275
rect 254 271 257 273
rect 259 271 261 273
rect 254 269 261 271
rect 234 262 239 269
rect 266 268 271 275
rect 287 271 291 275
rect 332 275 339 281
rect 314 273 321 275
rect 314 271 316 273
rect 318 271 321 273
rect 287 268 293 271
rect 266 262 273 268
rect 275 266 283 268
rect 275 264 278 266
rect 280 264 283 266
rect 275 262 283 264
rect 285 262 293 268
rect 295 268 300 271
rect 314 269 321 271
rect 295 266 302 268
rect 295 264 298 266
rect 300 264 302 266
rect 316 264 321 269
rect 323 264 328 275
rect 330 273 339 275
rect 366 275 371 282
rect 364 273 371 275
rect 330 264 341 273
rect 343 271 350 273
rect 343 269 346 271
rect 348 269 350 271
rect 364 271 366 273
rect 368 271 371 273
rect 364 269 371 271
rect 373 279 378 282
rect 373 277 381 279
rect 373 275 376 277
rect 378 275 381 277
rect 373 269 381 275
rect 383 276 388 279
rect 383 274 391 276
rect 383 272 386 274
rect 388 272 391 274
rect 383 269 391 272
rect 343 267 350 269
rect 343 264 348 267
rect 295 262 302 264
rect 386 262 391 269
rect 393 266 401 276
rect 393 264 396 266
rect 398 264 401 266
rect 393 262 401 264
rect 403 273 410 276
rect 416 275 421 282
rect 403 271 406 273
rect 408 271 410 273
rect 403 266 410 271
rect 414 273 421 275
rect 414 271 416 273
rect 418 271 421 273
rect 414 269 421 271
rect 403 264 406 266
rect 408 264 410 266
rect 403 262 410 264
rect 416 262 421 269
rect 423 262 428 282
rect 430 280 439 282
rect 430 278 433 280
rect 435 278 439 280
rect 430 268 439 278
rect 441 275 446 282
rect 456 275 461 282
rect 441 273 448 275
rect 441 271 444 273
rect 446 271 448 273
rect 441 268 448 271
rect 454 273 461 275
rect 454 271 456 273
rect 458 271 461 273
rect 454 268 461 271
rect 463 280 472 282
rect 463 278 467 280
rect 469 278 472 280
rect 463 268 472 278
rect 430 262 437 268
rect 465 262 472 268
rect 474 262 479 282
rect 481 275 486 282
rect 524 279 529 282
rect 514 276 519 279
rect 481 273 488 275
rect 481 271 484 273
rect 486 271 488 273
rect 481 269 488 271
rect 492 273 499 276
rect 492 271 494 273
rect 496 271 499 273
rect 481 262 486 269
rect 492 266 499 271
rect 492 264 494 266
rect 496 264 499 266
rect 492 262 499 264
rect 501 266 509 276
rect 501 264 504 266
rect 506 264 509 266
rect 501 262 509 264
rect 511 274 519 276
rect 511 272 514 274
rect 516 272 519 274
rect 511 269 519 272
rect 521 277 529 279
rect 521 275 524 277
rect 526 275 529 277
rect 521 269 529 275
rect 531 275 536 282
rect 543 279 549 281
rect 543 277 545 279
rect 547 277 549 279
rect 543 275 549 277
rect 562 279 568 281
rect 609 283 616 285
rect 609 281 612 283
rect 614 281 616 283
rect 562 277 564 279
rect 566 277 568 279
rect 562 275 568 277
rect 531 273 538 275
rect 531 271 534 273
rect 536 271 538 273
rect 531 269 538 271
rect 511 262 516 269
rect 543 268 548 275
rect 564 271 568 275
rect 609 275 616 281
rect 591 273 598 275
rect 591 271 593 273
rect 595 271 598 273
rect 564 268 570 271
rect 543 262 550 268
rect 552 266 560 268
rect 552 264 555 266
rect 557 264 560 266
rect 552 262 560 264
rect 562 262 570 268
rect 572 268 577 271
rect 591 269 598 271
rect 572 266 579 268
rect 572 264 575 266
rect 577 264 579 266
rect 593 264 598 269
rect 600 264 605 275
rect 607 273 616 275
rect 642 275 647 282
rect 640 273 647 275
rect 607 264 618 273
rect 620 271 627 273
rect 620 269 623 271
rect 625 269 627 271
rect 640 271 642 273
rect 644 271 647 273
rect 640 269 647 271
rect 649 279 654 282
rect 649 277 657 279
rect 649 275 652 277
rect 654 275 657 277
rect 649 269 657 275
rect 659 276 664 279
rect 659 274 667 276
rect 659 272 662 274
rect 664 272 667 274
rect 659 269 667 272
rect 620 267 627 269
rect 620 264 625 267
rect 572 262 579 264
rect 662 262 667 269
rect 669 266 677 276
rect 669 264 672 266
rect 674 264 677 266
rect 669 262 677 264
rect 679 273 686 276
rect 692 275 697 282
rect 679 271 682 273
rect 684 271 686 273
rect 679 266 686 271
rect 690 273 697 275
rect 690 271 692 273
rect 694 271 697 273
rect 690 269 697 271
rect 679 264 682 266
rect 684 264 686 266
rect 679 262 686 264
rect 692 262 697 269
rect 699 262 704 282
rect 706 280 715 282
rect 706 278 709 280
rect 711 278 715 280
rect 706 268 715 278
rect 717 275 722 282
rect 732 275 737 282
rect 717 273 724 275
rect 717 271 720 273
rect 722 271 724 273
rect 717 268 724 271
rect 730 273 737 275
rect 730 271 732 273
rect 734 271 737 273
rect 730 268 737 271
rect 739 280 748 282
rect 739 278 743 280
rect 745 278 748 280
rect 739 268 748 278
rect 706 262 713 268
rect 741 262 748 268
rect 750 262 755 282
rect 757 275 762 282
rect 800 279 805 282
rect 790 276 795 279
rect 757 273 764 275
rect 757 271 760 273
rect 762 271 764 273
rect 757 269 764 271
rect 768 273 775 276
rect 768 271 770 273
rect 772 271 775 273
rect 757 262 762 269
rect 768 266 775 271
rect 768 264 770 266
rect 772 264 775 266
rect 768 262 775 264
rect 777 266 785 276
rect 777 264 780 266
rect 782 264 785 266
rect 777 262 785 264
rect 787 274 795 276
rect 787 272 790 274
rect 792 272 795 274
rect 787 269 795 272
rect 797 277 805 279
rect 797 275 800 277
rect 802 275 805 277
rect 797 269 805 275
rect 807 275 812 282
rect 819 279 825 281
rect 819 277 821 279
rect 823 277 825 279
rect 819 275 825 277
rect 838 279 844 281
rect 885 283 892 285
rect 885 281 888 283
rect 890 281 892 283
rect 838 277 840 279
rect 842 277 844 279
rect 838 275 844 277
rect 807 273 814 275
rect 807 271 810 273
rect 812 271 814 273
rect 807 269 814 271
rect 787 262 792 269
rect 819 268 824 275
rect 840 271 844 275
rect 885 275 892 281
rect 867 273 874 275
rect 867 271 869 273
rect 871 271 874 273
rect 840 268 846 271
rect 819 262 826 268
rect 828 266 836 268
rect 828 264 831 266
rect 833 264 836 266
rect 828 262 836 264
rect 838 262 846 268
rect 848 268 853 271
rect 867 269 874 271
rect 848 266 855 268
rect 848 264 851 266
rect 853 264 855 266
rect 869 264 874 269
rect 876 264 881 275
rect 883 273 892 275
rect 919 275 924 282
rect 917 273 924 275
rect 883 264 894 273
rect 896 271 903 273
rect 896 269 899 271
rect 901 269 903 271
rect 917 271 919 273
rect 921 271 924 273
rect 917 269 924 271
rect 926 279 931 282
rect 926 277 934 279
rect 926 275 929 277
rect 931 275 934 277
rect 926 269 934 275
rect 936 276 941 279
rect 936 274 944 276
rect 936 272 939 274
rect 941 272 944 274
rect 936 269 944 272
rect 896 267 903 269
rect 896 264 901 267
rect 848 262 855 264
rect 939 262 944 269
rect 946 266 954 276
rect 946 264 949 266
rect 951 264 954 266
rect 946 262 954 264
rect 956 273 963 276
rect 969 275 974 282
rect 956 271 959 273
rect 961 271 963 273
rect 956 266 963 271
rect 967 273 974 275
rect 967 271 969 273
rect 971 271 974 273
rect 967 269 974 271
rect 956 264 959 266
rect 961 264 963 266
rect 956 262 963 264
rect 969 262 974 269
rect 976 262 981 282
rect 983 280 992 282
rect 983 278 986 280
rect 988 278 992 280
rect 983 268 992 278
rect 994 275 999 282
rect 1009 275 1014 282
rect 994 273 1001 275
rect 994 271 997 273
rect 999 271 1001 273
rect 994 268 1001 271
rect 1007 273 1014 275
rect 1007 271 1009 273
rect 1011 271 1014 273
rect 1007 268 1014 271
rect 1016 280 1025 282
rect 1016 278 1020 280
rect 1022 278 1025 280
rect 1016 268 1025 278
rect 983 262 990 268
rect 1018 262 1025 268
rect 1027 262 1032 282
rect 1034 275 1039 282
rect 1077 279 1082 282
rect 1067 276 1072 279
rect 1034 273 1041 275
rect 1034 271 1037 273
rect 1039 271 1041 273
rect 1034 269 1041 271
rect 1045 273 1052 276
rect 1045 271 1047 273
rect 1049 271 1052 273
rect 1034 262 1039 269
rect 1045 266 1052 271
rect 1045 264 1047 266
rect 1049 264 1052 266
rect 1045 262 1052 264
rect 1054 266 1062 276
rect 1054 264 1057 266
rect 1059 264 1062 266
rect 1054 262 1062 264
rect 1064 274 1072 276
rect 1064 272 1067 274
rect 1069 272 1072 274
rect 1064 269 1072 272
rect 1074 277 1082 279
rect 1074 275 1077 277
rect 1079 275 1082 277
rect 1074 269 1082 275
rect 1084 275 1089 282
rect 1096 279 1102 281
rect 1096 277 1098 279
rect 1100 277 1102 279
rect 1096 275 1102 277
rect 1115 279 1121 281
rect 1115 277 1117 279
rect 1119 277 1121 279
rect 1115 275 1121 277
rect 1084 273 1091 275
rect 1084 271 1087 273
rect 1089 271 1091 273
rect 1084 269 1091 271
rect 1064 262 1069 269
rect 1096 268 1101 275
rect 1117 271 1121 275
rect 1117 268 1123 271
rect 1096 262 1103 268
rect 1105 266 1113 268
rect 1105 264 1108 266
rect 1110 264 1113 266
rect 1105 262 1113 264
rect 1115 262 1123 268
rect 1125 268 1130 271
rect 1125 266 1132 268
rect 1125 264 1128 266
rect 1130 264 1132 266
rect 1125 262 1132 264
rect -283 168 -276 170
rect -283 166 -281 168
rect -279 166 -276 168
rect -283 164 -276 166
rect -281 161 -276 164
rect -274 165 -269 170
rect -274 161 -260 165
rect -269 160 -260 161
rect -269 158 -267 160
rect -265 158 -260 160
rect -269 156 -260 158
rect -258 163 -250 165
rect -258 161 -255 163
rect -253 161 -250 163
rect -258 156 -250 161
rect -248 161 -240 165
rect -248 159 -245 161
rect -243 159 -240 161
rect -248 156 -240 159
rect -245 153 -240 156
rect -238 153 -233 165
rect -231 153 -223 165
rect -193 163 -188 170
rect -215 161 -208 163
rect -215 159 -213 161
rect -211 159 -208 161
rect -215 157 -208 159
rect -229 151 -223 153
rect -229 149 -227 151
rect -225 149 -223 151
rect -213 150 -208 157
rect -206 157 -198 163
rect -206 155 -203 157
rect -201 155 -198 157
rect -206 153 -198 155
rect -196 160 -188 163
rect -196 158 -193 160
rect -191 158 -188 160
rect -196 156 -188 158
rect -186 168 -178 170
rect -186 166 -183 168
rect -181 166 -178 168
rect -186 156 -178 166
rect -176 168 -169 170
rect -176 166 -173 168
rect -171 166 -169 168
rect -176 161 -169 166
rect -163 163 -158 170
rect -176 159 -173 161
rect -171 159 -169 161
rect -176 156 -169 159
rect -165 161 -158 163
rect -165 159 -163 161
rect -161 159 -158 161
rect -165 157 -158 159
rect -196 153 -191 156
rect -206 150 -201 153
rect -229 147 -223 149
rect -163 150 -158 157
rect -156 150 -151 170
rect -149 164 -142 170
rect -114 164 -107 170
rect -149 154 -140 164
rect -149 152 -146 154
rect -144 152 -140 154
rect -149 150 -140 152
rect -138 161 -131 164
rect -138 159 -135 161
rect -133 159 -131 161
rect -138 157 -131 159
rect -125 161 -118 164
rect -125 159 -123 161
rect -121 159 -118 161
rect -125 157 -118 159
rect -138 150 -133 157
rect -123 150 -118 157
rect -116 154 -107 164
rect -116 152 -112 154
rect -110 152 -107 154
rect -116 150 -107 152
rect -105 150 -100 170
rect -98 163 -93 170
rect -87 168 -80 170
rect -87 166 -85 168
rect -83 166 -80 168
rect -98 161 -91 163
rect -98 159 -95 161
rect -93 159 -91 161
rect -98 157 -91 159
rect -87 161 -80 166
rect -87 159 -85 161
rect -83 159 -80 161
rect -98 150 -93 157
rect -87 156 -80 159
rect -78 168 -70 170
rect -78 166 -75 168
rect -73 166 -70 168
rect -78 156 -70 166
rect -68 163 -63 170
rect -36 164 -29 170
rect -27 168 -19 170
rect -27 166 -24 168
rect -22 166 -19 168
rect -27 164 -19 166
rect -17 164 -9 170
rect -68 160 -60 163
rect -68 158 -65 160
rect -63 158 -60 160
rect -68 156 -60 158
rect -65 153 -60 156
rect -58 157 -50 163
rect -58 155 -55 157
rect -53 155 -50 157
rect -58 153 -50 155
rect -55 150 -50 153
rect -48 161 -41 163
rect -48 159 -45 161
rect -43 159 -41 161
rect -48 157 -41 159
rect -36 157 -31 164
rect -15 161 -9 164
rect -7 168 0 170
rect -7 166 -4 168
rect -2 166 0 168
rect -7 164 0 166
rect -7 161 -2 164
rect 9 163 14 168
rect 7 161 14 163
rect -15 157 -11 161
rect -48 150 -43 157
rect -36 155 -30 157
rect -36 153 -34 155
rect -32 153 -30 155
rect -36 151 -30 153
rect -17 155 -11 157
rect 7 159 9 161
rect 11 159 14 161
rect 7 157 14 159
rect 16 157 21 168
rect 23 159 34 168
rect 36 165 41 168
rect 36 163 43 165
rect 49 163 54 168
rect 36 161 39 163
rect 41 161 43 163
rect 36 159 43 161
rect 47 161 54 163
rect 47 159 49 161
rect 51 159 54 161
rect 23 157 32 159
rect -17 153 -15 155
rect -13 153 -11 155
rect -17 151 -11 153
rect 25 151 32 157
rect 47 157 54 159
rect 56 157 61 168
rect 63 159 74 168
rect 76 165 81 168
rect 76 163 83 165
rect 109 163 114 170
rect 76 161 79 163
rect 81 161 83 163
rect 76 159 83 161
rect 87 161 94 163
rect 87 159 89 161
rect 91 159 94 161
rect 63 157 72 159
rect 25 149 28 151
rect 30 149 32 151
rect 25 147 32 149
rect 65 151 72 157
rect 87 157 94 159
rect 65 149 68 151
rect 70 149 72 151
rect 65 147 72 149
rect 89 150 94 157
rect 96 157 104 163
rect 96 155 99 157
rect 101 155 104 157
rect 96 153 104 155
rect 106 160 114 163
rect 106 158 109 160
rect 111 158 114 160
rect 106 156 114 158
rect 116 168 124 170
rect 116 166 119 168
rect 121 166 124 168
rect 116 156 124 166
rect 126 168 133 170
rect 126 166 129 168
rect 131 166 133 168
rect 126 161 133 166
rect 139 163 144 170
rect 126 159 129 161
rect 131 159 133 161
rect 126 156 133 159
rect 137 161 144 163
rect 137 159 139 161
rect 141 159 144 161
rect 137 157 144 159
rect 106 153 111 156
rect 96 150 101 153
rect 139 150 144 157
rect 146 150 151 170
rect 153 164 160 170
rect 188 164 195 170
rect 153 154 162 164
rect 153 152 156 154
rect 158 152 162 154
rect 153 150 162 152
rect 164 161 171 164
rect 164 159 167 161
rect 169 159 171 161
rect 164 157 171 159
rect 177 161 184 164
rect 177 159 179 161
rect 181 159 184 161
rect 177 157 184 159
rect 164 150 169 157
rect 179 150 184 157
rect 186 154 195 164
rect 186 152 190 154
rect 192 152 195 154
rect 186 150 195 152
rect 197 150 202 170
rect 204 163 209 170
rect 215 168 222 170
rect 215 166 217 168
rect 219 166 222 168
rect 204 161 211 163
rect 204 159 207 161
rect 209 159 211 161
rect 204 157 211 159
rect 215 161 222 166
rect 215 159 217 161
rect 219 159 222 161
rect 204 150 209 157
rect 215 156 222 159
rect 224 168 232 170
rect 224 166 227 168
rect 229 166 232 168
rect 224 156 232 166
rect 234 163 239 170
rect 266 164 273 170
rect 275 168 283 170
rect 275 166 278 168
rect 280 166 283 168
rect 275 164 283 166
rect 285 164 293 170
rect 234 160 242 163
rect 234 158 237 160
rect 239 158 242 160
rect 234 156 242 158
rect 237 153 242 156
rect 244 157 252 163
rect 244 155 247 157
rect 249 155 252 157
rect 244 153 252 155
rect 247 150 252 153
rect 254 161 261 163
rect 254 159 257 161
rect 259 159 261 161
rect 254 157 261 159
rect 266 157 271 164
rect 287 161 293 164
rect 295 168 302 170
rect 295 166 298 168
rect 300 166 302 168
rect 295 164 302 166
rect 295 161 300 164
rect 316 163 321 168
rect 314 161 321 163
rect 287 157 291 161
rect 254 150 259 157
rect 266 155 272 157
rect 266 153 268 155
rect 270 153 272 155
rect 266 151 272 153
rect 285 155 291 157
rect 314 159 316 161
rect 318 159 321 161
rect 314 157 321 159
rect 323 157 328 168
rect 330 159 341 168
rect 343 165 348 168
rect 343 163 350 165
rect 386 163 391 170
rect 343 161 346 163
rect 348 161 350 163
rect 343 159 350 161
rect 364 161 371 163
rect 364 159 366 161
rect 368 159 371 161
rect 330 157 339 159
rect 285 153 287 155
rect 289 153 291 155
rect 285 151 291 153
rect 332 151 339 157
rect 364 157 371 159
rect 332 149 335 151
rect 337 149 339 151
rect 332 147 339 149
rect 366 150 371 157
rect 373 157 381 163
rect 373 155 376 157
rect 378 155 381 157
rect 373 153 381 155
rect 383 160 391 163
rect 383 158 386 160
rect 388 158 391 160
rect 383 156 391 158
rect 393 168 401 170
rect 393 166 396 168
rect 398 166 401 168
rect 393 156 401 166
rect 403 168 410 170
rect 403 166 406 168
rect 408 166 410 168
rect 403 161 410 166
rect 416 163 421 170
rect 403 159 406 161
rect 408 159 410 161
rect 403 156 410 159
rect 414 161 421 163
rect 414 159 416 161
rect 418 159 421 161
rect 414 157 421 159
rect 383 153 388 156
rect 373 150 378 153
rect 416 150 421 157
rect 423 150 428 170
rect 430 164 437 170
rect 465 164 472 170
rect 430 154 439 164
rect 430 152 433 154
rect 435 152 439 154
rect 430 150 439 152
rect 441 161 448 164
rect 441 159 444 161
rect 446 159 448 161
rect 441 157 448 159
rect 454 161 461 164
rect 454 159 456 161
rect 458 159 461 161
rect 454 157 461 159
rect 441 150 446 157
rect 456 150 461 157
rect 463 154 472 164
rect 463 152 467 154
rect 469 152 472 154
rect 463 150 472 152
rect 474 150 479 170
rect 481 163 486 170
rect 492 168 499 170
rect 492 166 494 168
rect 496 166 499 168
rect 481 161 488 163
rect 481 159 484 161
rect 486 159 488 161
rect 481 157 488 159
rect 492 161 499 166
rect 492 159 494 161
rect 496 159 499 161
rect 481 150 486 157
rect 492 156 499 159
rect 501 168 509 170
rect 501 166 504 168
rect 506 166 509 168
rect 501 156 509 166
rect 511 163 516 170
rect 543 164 550 170
rect 552 168 560 170
rect 552 166 555 168
rect 557 166 560 168
rect 552 164 560 166
rect 562 164 570 170
rect 511 160 519 163
rect 511 158 514 160
rect 516 158 519 160
rect 511 156 519 158
rect 514 153 519 156
rect 521 157 529 163
rect 521 155 524 157
rect 526 155 529 157
rect 521 153 529 155
rect 524 150 529 153
rect 531 161 538 163
rect 531 159 534 161
rect 536 159 538 161
rect 531 157 538 159
rect 543 157 548 164
rect 564 161 570 164
rect 572 168 579 170
rect 572 166 575 168
rect 577 166 579 168
rect 572 164 579 166
rect 572 161 577 164
rect 593 163 598 168
rect 591 161 598 163
rect 564 157 568 161
rect 531 150 536 157
rect 543 155 549 157
rect 543 153 545 155
rect 547 153 549 155
rect 543 151 549 153
rect 562 155 568 157
rect 591 159 593 161
rect 595 159 598 161
rect 591 157 598 159
rect 600 157 605 168
rect 607 159 618 168
rect 620 165 625 168
rect 620 163 627 165
rect 662 163 667 170
rect 620 161 623 163
rect 625 161 627 163
rect 620 159 627 161
rect 640 161 647 163
rect 640 159 642 161
rect 644 159 647 161
rect 607 157 616 159
rect 562 153 564 155
rect 566 153 568 155
rect 562 151 568 153
rect 609 151 616 157
rect 640 157 647 159
rect 609 149 612 151
rect 614 149 616 151
rect 609 147 616 149
rect 642 150 647 157
rect 649 157 657 163
rect 649 155 652 157
rect 654 155 657 157
rect 649 153 657 155
rect 659 160 667 163
rect 659 158 662 160
rect 664 158 667 160
rect 659 156 667 158
rect 669 168 677 170
rect 669 166 672 168
rect 674 166 677 168
rect 669 156 677 166
rect 679 168 686 170
rect 679 166 682 168
rect 684 166 686 168
rect 679 161 686 166
rect 692 163 697 170
rect 679 159 682 161
rect 684 159 686 161
rect 679 156 686 159
rect 690 161 697 163
rect 690 159 692 161
rect 694 159 697 161
rect 690 157 697 159
rect 659 153 664 156
rect 649 150 654 153
rect 692 150 697 157
rect 699 150 704 170
rect 706 164 713 170
rect 741 164 748 170
rect 706 154 715 164
rect 706 152 709 154
rect 711 152 715 154
rect 706 150 715 152
rect 717 161 724 164
rect 717 159 720 161
rect 722 159 724 161
rect 717 157 724 159
rect 730 161 737 164
rect 730 159 732 161
rect 734 159 737 161
rect 730 157 737 159
rect 717 150 722 157
rect 732 150 737 157
rect 739 154 748 164
rect 739 152 743 154
rect 745 152 748 154
rect 739 150 748 152
rect 750 150 755 170
rect 757 163 762 170
rect 768 168 775 170
rect 768 166 770 168
rect 772 166 775 168
rect 757 161 764 163
rect 757 159 760 161
rect 762 159 764 161
rect 757 157 764 159
rect 768 161 775 166
rect 768 159 770 161
rect 772 159 775 161
rect 757 150 762 157
rect 768 156 775 159
rect 777 168 785 170
rect 777 166 780 168
rect 782 166 785 168
rect 777 156 785 166
rect 787 163 792 170
rect 819 164 826 170
rect 828 168 836 170
rect 828 166 831 168
rect 833 166 836 168
rect 828 164 836 166
rect 838 164 846 170
rect 787 160 795 163
rect 787 158 790 160
rect 792 158 795 160
rect 787 156 795 158
rect 790 153 795 156
rect 797 157 805 163
rect 797 155 800 157
rect 802 155 805 157
rect 797 153 805 155
rect 800 150 805 153
rect 807 161 814 163
rect 807 159 810 161
rect 812 159 814 161
rect 807 157 814 159
rect 819 157 824 164
rect 840 161 846 164
rect 848 168 855 170
rect 848 166 851 168
rect 853 166 855 168
rect 848 164 855 166
rect 848 161 853 164
rect 869 163 874 168
rect 867 161 874 163
rect 840 157 844 161
rect 807 150 812 157
rect 819 155 825 157
rect 819 153 821 155
rect 823 153 825 155
rect 819 151 825 153
rect 838 155 844 157
rect 867 159 869 161
rect 871 159 874 161
rect 867 157 874 159
rect 876 157 881 168
rect 883 159 894 168
rect 896 165 901 168
rect 896 163 903 165
rect 939 163 944 170
rect 896 161 899 163
rect 901 161 903 163
rect 896 159 903 161
rect 917 161 924 163
rect 917 159 919 161
rect 921 159 924 161
rect 883 157 892 159
rect 838 153 840 155
rect 842 153 844 155
rect 838 151 844 153
rect 885 151 892 157
rect 917 157 924 159
rect 885 149 888 151
rect 890 149 892 151
rect 885 147 892 149
rect 919 150 924 157
rect 926 157 934 163
rect 926 155 929 157
rect 931 155 934 157
rect 926 153 934 155
rect 936 160 944 163
rect 936 158 939 160
rect 941 158 944 160
rect 936 156 944 158
rect 946 168 954 170
rect 946 166 949 168
rect 951 166 954 168
rect 946 156 954 166
rect 956 168 963 170
rect 956 166 959 168
rect 961 166 963 168
rect 956 161 963 166
rect 969 163 974 170
rect 956 159 959 161
rect 961 159 963 161
rect 956 156 963 159
rect 967 161 974 163
rect 967 159 969 161
rect 971 159 974 161
rect 967 157 974 159
rect 936 153 941 156
rect 926 150 931 153
rect 969 150 974 157
rect 976 150 981 170
rect 983 164 990 170
rect 1018 164 1025 170
rect 983 154 992 164
rect 983 152 986 154
rect 988 152 992 154
rect 983 150 992 152
rect 994 161 1001 164
rect 994 159 997 161
rect 999 159 1001 161
rect 994 157 1001 159
rect 1007 161 1014 164
rect 1007 159 1009 161
rect 1011 159 1014 161
rect 1007 157 1014 159
rect 994 150 999 157
rect 1009 150 1014 157
rect 1016 154 1025 164
rect 1016 152 1020 154
rect 1022 152 1025 154
rect 1016 150 1025 152
rect 1027 150 1032 170
rect 1034 163 1039 170
rect 1045 168 1052 170
rect 1045 166 1047 168
rect 1049 166 1052 168
rect 1034 161 1041 163
rect 1034 159 1037 161
rect 1039 159 1041 161
rect 1034 157 1041 159
rect 1045 161 1052 166
rect 1045 159 1047 161
rect 1049 159 1052 161
rect 1034 150 1039 157
rect 1045 156 1052 159
rect 1054 168 1062 170
rect 1054 166 1057 168
rect 1059 166 1062 168
rect 1054 156 1062 166
rect 1064 163 1069 170
rect 1096 164 1103 170
rect 1105 168 1113 170
rect 1105 166 1108 168
rect 1110 166 1113 168
rect 1105 164 1113 166
rect 1115 164 1123 170
rect 1064 160 1072 163
rect 1064 158 1067 160
rect 1069 158 1072 160
rect 1064 156 1072 158
rect 1067 153 1072 156
rect 1074 157 1082 163
rect 1074 155 1077 157
rect 1079 155 1082 157
rect 1074 153 1082 155
rect 1077 150 1082 153
rect 1084 161 1091 163
rect 1084 159 1087 161
rect 1089 159 1091 161
rect 1084 157 1091 159
rect 1096 157 1101 164
rect 1117 161 1123 164
rect 1125 168 1132 170
rect 1125 166 1128 168
rect 1130 166 1132 168
rect 1125 164 1132 166
rect 1125 161 1130 164
rect 1117 157 1121 161
rect 1084 150 1089 157
rect 1096 155 1102 157
rect 1096 153 1098 155
rect 1100 153 1102 155
rect 1096 151 1102 153
rect 1115 155 1121 157
rect 1115 153 1117 155
rect 1119 153 1121 155
rect 1115 151 1121 153
rect -229 139 -223 141
rect -229 137 -227 139
rect -225 137 -223 139
rect -229 135 -223 137
rect -245 132 -240 135
rect -269 130 -260 132
rect -269 128 -267 130
rect -265 128 -260 130
rect -269 127 -260 128
rect -281 124 -276 127
rect -283 122 -276 124
rect -283 120 -281 122
rect -279 120 -276 122
rect -283 118 -276 120
rect -274 123 -260 127
rect -258 127 -250 132
rect -258 125 -255 127
rect -253 125 -250 127
rect -258 123 -250 125
rect -248 129 -240 132
rect -248 127 -245 129
rect -243 127 -240 129
rect -248 123 -240 127
rect -238 123 -233 135
rect -231 123 -223 135
rect -213 131 -208 138
rect -215 129 -208 131
rect -215 127 -213 129
rect -211 127 -208 129
rect -215 125 -208 127
rect -206 135 -201 138
rect -206 133 -198 135
rect -206 131 -203 133
rect -201 131 -198 133
rect -206 125 -198 131
rect -196 132 -191 135
rect -196 130 -188 132
rect -196 128 -193 130
rect -191 128 -188 130
rect -196 125 -188 128
rect -274 118 -269 123
rect -193 118 -188 125
rect -186 122 -178 132
rect -186 120 -183 122
rect -181 120 -178 122
rect -186 118 -178 120
rect -176 129 -169 132
rect -163 131 -158 138
rect -176 127 -173 129
rect -171 127 -169 129
rect -176 122 -169 127
rect -165 129 -158 131
rect -165 127 -163 129
rect -161 127 -158 129
rect -165 125 -158 127
rect -176 120 -173 122
rect -171 120 -169 122
rect -176 118 -169 120
rect -163 118 -158 125
rect -156 118 -151 138
rect -149 136 -140 138
rect -149 134 -146 136
rect -144 134 -140 136
rect -149 124 -140 134
rect -138 131 -133 138
rect -123 131 -118 138
rect -138 129 -131 131
rect -138 127 -135 129
rect -133 127 -131 129
rect -138 124 -131 127
rect -125 129 -118 131
rect -125 127 -123 129
rect -121 127 -118 129
rect -125 124 -118 127
rect -116 136 -107 138
rect -116 134 -112 136
rect -110 134 -107 136
rect -116 124 -107 134
rect -149 118 -142 124
rect -114 118 -107 124
rect -105 118 -100 138
rect -98 131 -93 138
rect -55 135 -50 138
rect -65 132 -60 135
rect -98 129 -91 131
rect -98 127 -95 129
rect -93 127 -91 129
rect -98 125 -91 127
rect -87 129 -80 132
rect -87 127 -85 129
rect -83 127 -80 129
rect -98 118 -93 125
rect -87 122 -80 127
rect -87 120 -85 122
rect -83 120 -80 122
rect -87 118 -80 120
rect -78 122 -70 132
rect -78 120 -75 122
rect -73 120 -70 122
rect -78 118 -70 120
rect -68 130 -60 132
rect -68 128 -65 130
rect -63 128 -60 130
rect -68 125 -60 128
rect -58 133 -50 135
rect -58 131 -55 133
rect -53 131 -50 133
rect -58 125 -50 131
rect -48 131 -43 138
rect -36 135 -30 137
rect -36 133 -34 135
rect -32 133 -30 135
rect -36 131 -30 133
rect -17 135 -11 137
rect 25 139 32 141
rect 25 137 28 139
rect 30 137 32 139
rect -17 133 -15 135
rect -13 133 -11 135
rect -17 131 -11 133
rect -48 129 -41 131
rect -48 127 -45 129
rect -43 127 -41 129
rect -48 125 -41 127
rect -68 118 -63 125
rect -36 124 -31 131
rect -15 127 -11 131
rect 25 131 32 137
rect 65 139 72 141
rect 65 137 68 139
rect 70 137 72 139
rect 7 129 14 131
rect 7 127 9 129
rect 11 127 14 129
rect -15 124 -9 127
rect -36 118 -29 124
rect -27 122 -19 124
rect -27 120 -24 122
rect -22 120 -19 122
rect -27 118 -19 120
rect -17 118 -9 124
rect -7 124 -2 127
rect 7 125 14 127
rect -7 122 0 124
rect -7 120 -4 122
rect -2 120 0 122
rect 9 120 14 125
rect 16 120 21 131
rect 23 129 32 131
rect 65 131 72 137
rect 47 129 54 131
rect 23 120 34 129
rect 36 127 43 129
rect 36 125 39 127
rect 41 125 43 127
rect 47 127 49 129
rect 51 127 54 129
rect 47 125 54 127
rect 36 123 43 125
rect 36 120 41 123
rect 49 120 54 125
rect 56 120 61 131
rect 63 129 72 131
rect 89 131 94 138
rect 87 129 94 131
rect 63 120 74 129
rect 76 127 83 129
rect 76 125 79 127
rect 81 125 83 127
rect 87 127 89 129
rect 91 127 94 129
rect 87 125 94 127
rect 96 135 101 138
rect 96 133 104 135
rect 96 131 99 133
rect 101 131 104 133
rect 96 125 104 131
rect 106 132 111 135
rect 106 130 114 132
rect 106 128 109 130
rect 111 128 114 130
rect 106 125 114 128
rect 76 123 83 125
rect 76 120 81 123
rect -7 118 0 120
rect 109 118 114 125
rect 116 122 124 132
rect 116 120 119 122
rect 121 120 124 122
rect 116 118 124 120
rect 126 129 133 132
rect 139 131 144 138
rect 126 127 129 129
rect 131 127 133 129
rect 126 122 133 127
rect 137 129 144 131
rect 137 127 139 129
rect 141 127 144 129
rect 137 125 144 127
rect 126 120 129 122
rect 131 120 133 122
rect 126 118 133 120
rect 139 118 144 125
rect 146 118 151 138
rect 153 136 162 138
rect 153 134 156 136
rect 158 134 162 136
rect 153 124 162 134
rect 164 131 169 138
rect 179 131 184 138
rect 164 129 171 131
rect 164 127 167 129
rect 169 127 171 129
rect 164 124 171 127
rect 177 129 184 131
rect 177 127 179 129
rect 181 127 184 129
rect 177 124 184 127
rect 186 136 195 138
rect 186 134 190 136
rect 192 134 195 136
rect 186 124 195 134
rect 153 118 160 124
rect 188 118 195 124
rect 197 118 202 138
rect 204 131 209 138
rect 247 135 252 138
rect 237 132 242 135
rect 204 129 211 131
rect 204 127 207 129
rect 209 127 211 129
rect 204 125 211 127
rect 215 129 222 132
rect 215 127 217 129
rect 219 127 222 129
rect 204 118 209 125
rect 215 122 222 127
rect 215 120 217 122
rect 219 120 222 122
rect 215 118 222 120
rect 224 122 232 132
rect 224 120 227 122
rect 229 120 232 122
rect 224 118 232 120
rect 234 130 242 132
rect 234 128 237 130
rect 239 128 242 130
rect 234 125 242 128
rect 244 133 252 135
rect 244 131 247 133
rect 249 131 252 133
rect 244 125 252 131
rect 254 131 259 138
rect 266 135 272 137
rect 266 133 268 135
rect 270 133 272 135
rect 266 131 272 133
rect 285 135 291 137
rect 332 139 339 141
rect 332 137 335 139
rect 337 137 339 139
rect 285 133 287 135
rect 289 133 291 135
rect 285 131 291 133
rect 254 129 261 131
rect 254 127 257 129
rect 259 127 261 129
rect 254 125 261 127
rect 234 118 239 125
rect 266 124 271 131
rect 287 127 291 131
rect 332 131 339 137
rect 314 129 321 131
rect 314 127 316 129
rect 318 127 321 129
rect 287 124 293 127
rect 266 118 273 124
rect 275 122 283 124
rect 275 120 278 122
rect 280 120 283 122
rect 275 118 283 120
rect 285 118 293 124
rect 295 124 300 127
rect 314 125 321 127
rect 295 122 302 124
rect 295 120 298 122
rect 300 120 302 122
rect 316 120 321 125
rect 323 120 328 131
rect 330 129 339 131
rect 366 131 371 138
rect 364 129 371 131
rect 330 120 341 129
rect 343 127 350 129
rect 343 125 346 127
rect 348 125 350 127
rect 364 127 366 129
rect 368 127 371 129
rect 364 125 371 127
rect 373 135 378 138
rect 373 133 381 135
rect 373 131 376 133
rect 378 131 381 133
rect 373 125 381 131
rect 383 132 388 135
rect 383 130 391 132
rect 383 128 386 130
rect 388 128 391 130
rect 383 125 391 128
rect 343 123 350 125
rect 343 120 348 123
rect 295 118 302 120
rect 386 118 391 125
rect 393 122 401 132
rect 393 120 396 122
rect 398 120 401 122
rect 393 118 401 120
rect 403 129 410 132
rect 416 131 421 138
rect 403 127 406 129
rect 408 127 410 129
rect 403 122 410 127
rect 414 129 421 131
rect 414 127 416 129
rect 418 127 421 129
rect 414 125 421 127
rect 403 120 406 122
rect 408 120 410 122
rect 403 118 410 120
rect 416 118 421 125
rect 423 118 428 138
rect 430 136 439 138
rect 430 134 433 136
rect 435 134 439 136
rect 430 124 439 134
rect 441 131 446 138
rect 456 131 461 138
rect 441 129 448 131
rect 441 127 444 129
rect 446 127 448 129
rect 441 124 448 127
rect 454 129 461 131
rect 454 127 456 129
rect 458 127 461 129
rect 454 124 461 127
rect 463 136 472 138
rect 463 134 467 136
rect 469 134 472 136
rect 463 124 472 134
rect 430 118 437 124
rect 465 118 472 124
rect 474 118 479 138
rect 481 131 486 138
rect 524 135 529 138
rect 514 132 519 135
rect 481 129 488 131
rect 481 127 484 129
rect 486 127 488 129
rect 481 125 488 127
rect 492 129 499 132
rect 492 127 494 129
rect 496 127 499 129
rect 481 118 486 125
rect 492 122 499 127
rect 492 120 494 122
rect 496 120 499 122
rect 492 118 499 120
rect 501 122 509 132
rect 501 120 504 122
rect 506 120 509 122
rect 501 118 509 120
rect 511 130 519 132
rect 511 128 514 130
rect 516 128 519 130
rect 511 125 519 128
rect 521 133 529 135
rect 521 131 524 133
rect 526 131 529 133
rect 521 125 529 131
rect 531 131 536 138
rect 543 135 549 137
rect 543 133 545 135
rect 547 133 549 135
rect 543 131 549 133
rect 562 135 568 137
rect 609 139 616 141
rect 609 137 612 139
rect 614 137 616 139
rect 562 133 564 135
rect 566 133 568 135
rect 562 131 568 133
rect 531 129 538 131
rect 531 127 534 129
rect 536 127 538 129
rect 531 125 538 127
rect 511 118 516 125
rect 543 124 548 131
rect 564 127 568 131
rect 609 131 616 137
rect 591 129 598 131
rect 591 127 593 129
rect 595 127 598 129
rect 564 124 570 127
rect 543 118 550 124
rect 552 122 560 124
rect 552 120 555 122
rect 557 120 560 122
rect 552 118 560 120
rect 562 118 570 124
rect 572 124 577 127
rect 591 125 598 127
rect 572 122 579 124
rect 572 120 575 122
rect 577 120 579 122
rect 593 120 598 125
rect 600 120 605 131
rect 607 129 616 131
rect 642 131 647 138
rect 640 129 647 131
rect 607 120 618 129
rect 620 127 627 129
rect 620 125 623 127
rect 625 125 627 127
rect 640 127 642 129
rect 644 127 647 129
rect 640 125 647 127
rect 649 135 654 138
rect 649 133 657 135
rect 649 131 652 133
rect 654 131 657 133
rect 649 125 657 131
rect 659 132 664 135
rect 659 130 667 132
rect 659 128 662 130
rect 664 128 667 130
rect 659 125 667 128
rect 620 123 627 125
rect 620 120 625 123
rect 572 118 579 120
rect 662 118 667 125
rect 669 122 677 132
rect 669 120 672 122
rect 674 120 677 122
rect 669 118 677 120
rect 679 129 686 132
rect 692 131 697 138
rect 679 127 682 129
rect 684 127 686 129
rect 679 122 686 127
rect 690 129 697 131
rect 690 127 692 129
rect 694 127 697 129
rect 690 125 697 127
rect 679 120 682 122
rect 684 120 686 122
rect 679 118 686 120
rect 692 118 697 125
rect 699 118 704 138
rect 706 136 715 138
rect 706 134 709 136
rect 711 134 715 136
rect 706 124 715 134
rect 717 131 722 138
rect 732 131 737 138
rect 717 129 724 131
rect 717 127 720 129
rect 722 127 724 129
rect 717 124 724 127
rect 730 129 737 131
rect 730 127 732 129
rect 734 127 737 129
rect 730 124 737 127
rect 739 136 748 138
rect 739 134 743 136
rect 745 134 748 136
rect 739 124 748 134
rect 706 118 713 124
rect 741 118 748 124
rect 750 118 755 138
rect 757 131 762 138
rect 800 135 805 138
rect 790 132 795 135
rect 757 129 764 131
rect 757 127 760 129
rect 762 127 764 129
rect 757 125 764 127
rect 768 129 775 132
rect 768 127 770 129
rect 772 127 775 129
rect 757 118 762 125
rect 768 122 775 127
rect 768 120 770 122
rect 772 120 775 122
rect 768 118 775 120
rect 777 122 785 132
rect 777 120 780 122
rect 782 120 785 122
rect 777 118 785 120
rect 787 130 795 132
rect 787 128 790 130
rect 792 128 795 130
rect 787 125 795 128
rect 797 133 805 135
rect 797 131 800 133
rect 802 131 805 133
rect 797 125 805 131
rect 807 131 812 138
rect 819 135 825 137
rect 819 133 821 135
rect 823 133 825 135
rect 819 131 825 133
rect 838 135 844 137
rect 885 139 892 141
rect 885 137 888 139
rect 890 137 892 139
rect 838 133 840 135
rect 842 133 844 135
rect 838 131 844 133
rect 807 129 814 131
rect 807 127 810 129
rect 812 127 814 129
rect 807 125 814 127
rect 787 118 792 125
rect 819 124 824 131
rect 840 127 844 131
rect 885 131 892 137
rect 867 129 874 131
rect 867 127 869 129
rect 871 127 874 129
rect 840 124 846 127
rect 819 118 826 124
rect 828 122 836 124
rect 828 120 831 122
rect 833 120 836 122
rect 828 118 836 120
rect 838 118 846 124
rect 848 124 853 127
rect 867 125 874 127
rect 848 122 855 124
rect 848 120 851 122
rect 853 120 855 122
rect 869 120 874 125
rect 876 120 881 131
rect 883 129 892 131
rect 919 131 924 138
rect 917 129 924 131
rect 883 120 894 129
rect 896 127 903 129
rect 896 125 899 127
rect 901 125 903 127
rect 917 127 919 129
rect 921 127 924 129
rect 917 125 924 127
rect 926 135 931 138
rect 926 133 934 135
rect 926 131 929 133
rect 931 131 934 133
rect 926 125 934 131
rect 936 132 941 135
rect 936 130 944 132
rect 936 128 939 130
rect 941 128 944 130
rect 936 125 944 128
rect 896 123 903 125
rect 896 120 901 123
rect 848 118 855 120
rect 939 118 944 125
rect 946 122 954 132
rect 946 120 949 122
rect 951 120 954 122
rect 946 118 954 120
rect 956 129 963 132
rect 969 131 974 138
rect 956 127 959 129
rect 961 127 963 129
rect 956 122 963 127
rect 967 129 974 131
rect 967 127 969 129
rect 971 127 974 129
rect 967 125 974 127
rect 956 120 959 122
rect 961 120 963 122
rect 956 118 963 120
rect 969 118 974 125
rect 976 118 981 138
rect 983 136 992 138
rect 983 134 986 136
rect 988 134 992 136
rect 983 124 992 134
rect 994 131 999 138
rect 1009 131 1014 138
rect 994 129 1001 131
rect 994 127 997 129
rect 999 127 1001 129
rect 994 124 1001 127
rect 1007 129 1014 131
rect 1007 127 1009 129
rect 1011 127 1014 129
rect 1007 124 1014 127
rect 1016 136 1025 138
rect 1016 134 1020 136
rect 1022 134 1025 136
rect 1016 124 1025 134
rect 983 118 990 124
rect 1018 118 1025 124
rect 1027 118 1032 138
rect 1034 131 1039 138
rect 1077 135 1082 138
rect 1067 132 1072 135
rect 1034 129 1041 131
rect 1034 127 1037 129
rect 1039 127 1041 129
rect 1034 125 1041 127
rect 1045 129 1052 132
rect 1045 127 1047 129
rect 1049 127 1052 129
rect 1034 118 1039 125
rect 1045 122 1052 127
rect 1045 120 1047 122
rect 1049 120 1052 122
rect 1045 118 1052 120
rect 1054 122 1062 132
rect 1054 120 1057 122
rect 1059 120 1062 122
rect 1054 118 1062 120
rect 1064 130 1072 132
rect 1064 128 1067 130
rect 1069 128 1072 130
rect 1064 125 1072 128
rect 1074 133 1082 135
rect 1074 131 1077 133
rect 1079 131 1082 133
rect 1074 125 1082 131
rect 1084 131 1089 138
rect 1096 135 1102 137
rect 1096 133 1098 135
rect 1100 133 1102 135
rect 1096 131 1102 133
rect 1115 135 1121 137
rect 1115 133 1117 135
rect 1119 133 1121 135
rect 1115 131 1121 133
rect 1084 129 1091 131
rect 1084 127 1087 129
rect 1089 127 1091 129
rect 1084 125 1091 127
rect 1064 118 1069 125
rect 1096 124 1101 131
rect 1117 127 1121 131
rect 1117 124 1123 127
rect 1096 118 1103 124
rect 1105 122 1113 124
rect 1105 120 1108 122
rect 1110 120 1113 122
rect 1105 118 1113 120
rect 1115 118 1123 124
rect 1125 124 1130 127
rect 1125 122 1132 124
rect 1125 120 1128 122
rect 1130 120 1132 122
rect 1125 118 1132 120
rect -283 24 -276 26
rect -283 22 -281 24
rect -279 22 -276 24
rect -283 20 -276 22
rect -281 17 -276 20
rect -274 21 -269 26
rect -274 17 -260 21
rect -269 16 -260 17
rect -269 14 -267 16
rect -265 14 -260 16
rect -269 12 -260 14
rect -258 19 -250 21
rect -258 17 -255 19
rect -253 17 -250 19
rect -258 12 -250 17
rect -248 17 -240 21
rect -248 15 -245 17
rect -243 15 -240 17
rect -248 12 -240 15
rect -245 9 -240 12
rect -238 9 -233 21
rect -231 9 -223 21
rect -193 19 -188 26
rect -215 17 -208 19
rect -215 15 -213 17
rect -211 15 -208 17
rect -215 13 -208 15
rect -229 7 -223 9
rect -229 5 -227 7
rect -225 5 -223 7
rect -213 6 -208 13
rect -206 13 -198 19
rect -206 11 -203 13
rect -201 11 -198 13
rect -206 9 -198 11
rect -196 16 -188 19
rect -196 14 -193 16
rect -191 14 -188 16
rect -196 12 -188 14
rect -186 24 -178 26
rect -186 22 -183 24
rect -181 22 -178 24
rect -186 12 -178 22
rect -176 24 -169 26
rect -176 22 -173 24
rect -171 22 -169 24
rect -176 17 -169 22
rect -163 19 -158 26
rect -176 15 -173 17
rect -171 15 -169 17
rect -176 12 -169 15
rect -165 17 -158 19
rect -165 15 -163 17
rect -161 15 -158 17
rect -165 13 -158 15
rect -196 9 -191 12
rect -206 6 -201 9
rect -229 3 -223 5
rect -163 6 -158 13
rect -156 6 -151 26
rect -149 20 -142 26
rect -114 20 -107 26
rect -149 10 -140 20
rect -149 8 -146 10
rect -144 8 -140 10
rect -149 6 -140 8
rect -138 17 -131 20
rect -138 15 -135 17
rect -133 15 -131 17
rect -138 13 -131 15
rect -125 17 -118 20
rect -125 15 -123 17
rect -121 15 -118 17
rect -125 13 -118 15
rect -138 6 -133 13
rect -123 6 -118 13
rect -116 10 -107 20
rect -116 8 -112 10
rect -110 8 -107 10
rect -116 6 -107 8
rect -105 6 -100 26
rect -98 19 -93 26
rect -87 24 -80 26
rect -87 22 -85 24
rect -83 22 -80 24
rect -98 17 -91 19
rect -98 15 -95 17
rect -93 15 -91 17
rect -98 13 -91 15
rect -87 17 -80 22
rect -87 15 -85 17
rect -83 15 -80 17
rect -98 6 -93 13
rect -87 12 -80 15
rect -78 24 -70 26
rect -78 22 -75 24
rect -73 22 -70 24
rect -78 12 -70 22
rect -68 19 -63 26
rect -36 20 -29 26
rect -27 24 -19 26
rect -27 22 -24 24
rect -22 22 -19 24
rect -27 20 -19 22
rect -17 20 -9 26
rect -68 16 -60 19
rect -68 14 -65 16
rect -63 14 -60 16
rect -68 12 -60 14
rect -65 9 -60 12
rect -58 13 -50 19
rect -58 11 -55 13
rect -53 11 -50 13
rect -58 9 -50 11
rect -55 6 -50 9
rect -48 17 -41 19
rect -48 15 -45 17
rect -43 15 -41 17
rect -48 13 -41 15
rect -36 13 -31 20
rect -15 17 -9 20
rect -7 24 0 26
rect -7 22 -4 24
rect -2 22 0 24
rect -7 20 0 22
rect -7 17 -2 20
rect 9 19 14 24
rect 7 17 14 19
rect -15 13 -11 17
rect -48 6 -43 13
rect -36 11 -30 13
rect -36 9 -34 11
rect -32 9 -30 11
rect -36 7 -30 9
rect -17 11 -11 13
rect 7 15 9 17
rect 11 15 14 17
rect 7 13 14 15
rect 16 13 21 24
rect 23 15 34 24
rect 36 21 41 24
rect 36 19 43 21
rect 49 19 54 24
rect 36 17 39 19
rect 41 17 43 19
rect 36 15 43 17
rect 47 17 54 19
rect 47 15 49 17
rect 51 15 54 17
rect 23 13 32 15
rect -17 9 -15 11
rect -13 9 -11 11
rect -17 7 -11 9
rect 25 7 32 13
rect 47 13 54 15
rect 56 13 61 24
rect 63 15 74 24
rect 76 21 81 24
rect 76 19 83 21
rect 109 19 114 26
rect 76 17 79 19
rect 81 17 83 19
rect 76 15 83 17
rect 87 17 94 19
rect 87 15 89 17
rect 91 15 94 17
rect 63 13 72 15
rect 25 5 28 7
rect 30 5 32 7
rect 25 3 32 5
rect 65 7 72 13
rect 87 13 94 15
rect 65 5 68 7
rect 70 5 72 7
rect 65 3 72 5
rect 89 6 94 13
rect 96 13 104 19
rect 96 11 99 13
rect 101 11 104 13
rect 96 9 104 11
rect 106 16 114 19
rect 106 14 109 16
rect 111 14 114 16
rect 106 12 114 14
rect 116 24 124 26
rect 116 22 119 24
rect 121 22 124 24
rect 116 12 124 22
rect 126 24 133 26
rect 126 22 129 24
rect 131 22 133 24
rect 126 17 133 22
rect 139 19 144 26
rect 126 15 129 17
rect 131 15 133 17
rect 126 12 133 15
rect 137 17 144 19
rect 137 15 139 17
rect 141 15 144 17
rect 137 13 144 15
rect 106 9 111 12
rect 96 6 101 9
rect 139 6 144 13
rect 146 6 151 26
rect 153 20 160 26
rect 188 20 195 26
rect 153 10 162 20
rect 153 8 156 10
rect 158 8 162 10
rect 153 6 162 8
rect 164 17 171 20
rect 164 15 167 17
rect 169 15 171 17
rect 164 13 171 15
rect 177 17 184 20
rect 177 15 179 17
rect 181 15 184 17
rect 177 13 184 15
rect 164 6 169 13
rect 179 6 184 13
rect 186 10 195 20
rect 186 8 190 10
rect 192 8 195 10
rect 186 6 195 8
rect 197 6 202 26
rect 204 19 209 26
rect 215 24 222 26
rect 215 22 217 24
rect 219 22 222 24
rect 204 17 211 19
rect 204 15 207 17
rect 209 15 211 17
rect 204 13 211 15
rect 215 17 222 22
rect 215 15 217 17
rect 219 15 222 17
rect 204 6 209 13
rect 215 12 222 15
rect 224 24 232 26
rect 224 22 227 24
rect 229 22 232 24
rect 224 12 232 22
rect 234 19 239 26
rect 266 20 273 26
rect 275 24 283 26
rect 275 22 278 24
rect 280 22 283 24
rect 275 20 283 22
rect 285 20 293 26
rect 234 16 242 19
rect 234 14 237 16
rect 239 14 242 16
rect 234 12 242 14
rect 237 9 242 12
rect 244 13 252 19
rect 244 11 247 13
rect 249 11 252 13
rect 244 9 252 11
rect 247 6 252 9
rect 254 17 261 19
rect 254 15 257 17
rect 259 15 261 17
rect 254 13 261 15
rect 266 13 271 20
rect 287 17 293 20
rect 295 24 302 26
rect 295 22 298 24
rect 300 22 302 24
rect 295 20 302 22
rect 295 17 300 20
rect 316 19 321 24
rect 314 17 321 19
rect 287 13 291 17
rect 254 6 259 13
rect 266 11 272 13
rect 266 9 268 11
rect 270 9 272 11
rect 266 7 272 9
rect 285 11 291 13
rect 314 15 316 17
rect 318 15 321 17
rect 314 13 321 15
rect 323 13 328 24
rect 330 15 341 24
rect 343 21 348 24
rect 343 19 350 21
rect 386 19 391 26
rect 343 17 346 19
rect 348 17 350 19
rect 343 15 350 17
rect 364 17 371 19
rect 364 15 366 17
rect 368 15 371 17
rect 330 13 339 15
rect 285 9 287 11
rect 289 9 291 11
rect 285 7 291 9
rect 332 7 339 13
rect 364 13 371 15
rect 332 5 335 7
rect 337 5 339 7
rect 332 3 339 5
rect 366 6 371 13
rect 373 13 381 19
rect 373 11 376 13
rect 378 11 381 13
rect 373 9 381 11
rect 383 16 391 19
rect 383 14 386 16
rect 388 14 391 16
rect 383 12 391 14
rect 393 24 401 26
rect 393 22 396 24
rect 398 22 401 24
rect 393 12 401 22
rect 403 24 410 26
rect 403 22 406 24
rect 408 22 410 24
rect 403 17 410 22
rect 416 19 421 26
rect 403 15 406 17
rect 408 15 410 17
rect 403 12 410 15
rect 414 17 421 19
rect 414 15 416 17
rect 418 15 421 17
rect 414 13 421 15
rect 383 9 388 12
rect 373 6 378 9
rect 416 6 421 13
rect 423 6 428 26
rect 430 20 437 26
rect 465 20 472 26
rect 430 10 439 20
rect 430 8 433 10
rect 435 8 439 10
rect 430 6 439 8
rect 441 17 448 20
rect 441 15 444 17
rect 446 15 448 17
rect 441 13 448 15
rect 454 17 461 20
rect 454 15 456 17
rect 458 15 461 17
rect 454 13 461 15
rect 441 6 446 13
rect 456 6 461 13
rect 463 10 472 20
rect 463 8 467 10
rect 469 8 472 10
rect 463 6 472 8
rect 474 6 479 26
rect 481 19 486 26
rect 492 24 499 26
rect 492 22 494 24
rect 496 22 499 24
rect 481 17 488 19
rect 481 15 484 17
rect 486 15 488 17
rect 481 13 488 15
rect 492 17 499 22
rect 492 15 494 17
rect 496 15 499 17
rect 481 6 486 13
rect 492 12 499 15
rect 501 24 509 26
rect 501 22 504 24
rect 506 22 509 24
rect 501 12 509 22
rect 511 19 516 26
rect 543 20 550 26
rect 552 24 560 26
rect 552 22 555 24
rect 557 22 560 24
rect 552 20 560 22
rect 562 20 570 26
rect 511 16 519 19
rect 511 14 514 16
rect 516 14 519 16
rect 511 12 519 14
rect 514 9 519 12
rect 521 13 529 19
rect 521 11 524 13
rect 526 11 529 13
rect 521 9 529 11
rect 524 6 529 9
rect 531 17 538 19
rect 531 15 534 17
rect 536 15 538 17
rect 531 13 538 15
rect 543 13 548 20
rect 564 17 570 20
rect 572 24 579 26
rect 572 22 575 24
rect 577 22 579 24
rect 572 20 579 22
rect 572 17 577 20
rect 593 19 598 24
rect 591 17 598 19
rect 564 13 568 17
rect 531 6 536 13
rect 543 11 549 13
rect 543 9 545 11
rect 547 9 549 11
rect 543 7 549 9
rect 562 11 568 13
rect 591 15 593 17
rect 595 15 598 17
rect 591 13 598 15
rect 600 13 605 24
rect 607 15 618 24
rect 620 21 625 24
rect 620 19 627 21
rect 662 19 667 26
rect 620 17 623 19
rect 625 17 627 19
rect 620 15 627 17
rect 640 17 647 19
rect 640 15 642 17
rect 644 15 647 17
rect 607 13 616 15
rect 562 9 564 11
rect 566 9 568 11
rect 562 7 568 9
rect 609 7 616 13
rect 640 13 647 15
rect 609 5 612 7
rect 614 5 616 7
rect 609 3 616 5
rect 642 6 647 13
rect 649 13 657 19
rect 649 11 652 13
rect 654 11 657 13
rect 649 9 657 11
rect 659 16 667 19
rect 659 14 662 16
rect 664 14 667 16
rect 659 12 667 14
rect 669 24 677 26
rect 669 22 672 24
rect 674 22 677 24
rect 669 12 677 22
rect 679 24 686 26
rect 679 22 682 24
rect 684 22 686 24
rect 679 17 686 22
rect 692 19 697 26
rect 679 15 682 17
rect 684 15 686 17
rect 679 12 686 15
rect 690 17 697 19
rect 690 15 692 17
rect 694 15 697 17
rect 690 13 697 15
rect 659 9 664 12
rect 649 6 654 9
rect 692 6 697 13
rect 699 6 704 26
rect 706 20 713 26
rect 741 20 748 26
rect 706 10 715 20
rect 706 8 709 10
rect 711 8 715 10
rect 706 6 715 8
rect 717 17 724 20
rect 717 15 720 17
rect 722 15 724 17
rect 717 13 724 15
rect 730 17 737 20
rect 730 15 732 17
rect 734 15 737 17
rect 730 13 737 15
rect 717 6 722 13
rect 732 6 737 13
rect 739 10 748 20
rect 739 8 743 10
rect 745 8 748 10
rect 739 6 748 8
rect 750 6 755 26
rect 757 19 762 26
rect 768 24 775 26
rect 768 22 770 24
rect 772 22 775 24
rect 757 17 764 19
rect 757 15 760 17
rect 762 15 764 17
rect 757 13 764 15
rect 768 17 775 22
rect 768 15 770 17
rect 772 15 775 17
rect 757 6 762 13
rect 768 12 775 15
rect 777 24 785 26
rect 777 22 780 24
rect 782 22 785 24
rect 777 12 785 22
rect 787 19 792 26
rect 819 20 826 26
rect 828 24 836 26
rect 828 22 831 24
rect 833 22 836 24
rect 828 20 836 22
rect 838 20 846 26
rect 787 16 795 19
rect 787 14 790 16
rect 792 14 795 16
rect 787 12 795 14
rect 790 9 795 12
rect 797 13 805 19
rect 797 11 800 13
rect 802 11 805 13
rect 797 9 805 11
rect 800 6 805 9
rect 807 17 814 19
rect 807 15 810 17
rect 812 15 814 17
rect 807 13 814 15
rect 819 13 824 20
rect 840 17 846 20
rect 848 24 855 26
rect 848 22 851 24
rect 853 22 855 24
rect 848 20 855 22
rect 848 17 853 20
rect 869 19 874 24
rect 867 17 874 19
rect 840 13 844 17
rect 807 6 812 13
rect 819 11 825 13
rect 819 9 821 11
rect 823 9 825 11
rect 819 7 825 9
rect 838 11 844 13
rect 867 15 869 17
rect 871 15 874 17
rect 867 13 874 15
rect 876 13 881 24
rect 883 15 894 24
rect 896 21 901 24
rect 896 19 903 21
rect 939 19 944 26
rect 896 17 899 19
rect 901 17 903 19
rect 896 15 903 17
rect 917 17 924 19
rect 917 15 919 17
rect 921 15 924 17
rect 883 13 892 15
rect 838 9 840 11
rect 842 9 844 11
rect 838 7 844 9
rect 885 7 892 13
rect 917 13 924 15
rect 885 5 888 7
rect 890 5 892 7
rect 885 3 892 5
rect 919 6 924 13
rect 926 13 934 19
rect 926 11 929 13
rect 931 11 934 13
rect 926 9 934 11
rect 936 16 944 19
rect 936 14 939 16
rect 941 14 944 16
rect 936 12 944 14
rect 946 24 954 26
rect 946 22 949 24
rect 951 22 954 24
rect 946 12 954 22
rect 956 24 963 26
rect 956 22 959 24
rect 961 22 963 24
rect 956 17 963 22
rect 969 19 974 26
rect 956 15 959 17
rect 961 15 963 17
rect 956 12 963 15
rect 967 17 974 19
rect 967 15 969 17
rect 971 15 974 17
rect 967 13 974 15
rect 936 9 941 12
rect 926 6 931 9
rect 969 6 974 13
rect 976 6 981 26
rect 983 20 990 26
rect 1018 20 1025 26
rect 983 10 992 20
rect 983 8 986 10
rect 988 8 992 10
rect 983 6 992 8
rect 994 17 1001 20
rect 994 15 997 17
rect 999 15 1001 17
rect 994 13 1001 15
rect 1007 17 1014 20
rect 1007 15 1009 17
rect 1011 15 1014 17
rect 1007 13 1014 15
rect 994 6 999 13
rect 1009 6 1014 13
rect 1016 10 1025 20
rect 1016 8 1020 10
rect 1022 8 1025 10
rect 1016 6 1025 8
rect 1027 6 1032 26
rect 1034 19 1039 26
rect 1045 24 1052 26
rect 1045 22 1047 24
rect 1049 22 1052 24
rect 1034 17 1041 19
rect 1034 15 1037 17
rect 1039 15 1041 17
rect 1034 13 1041 15
rect 1045 17 1052 22
rect 1045 15 1047 17
rect 1049 15 1052 17
rect 1034 6 1039 13
rect 1045 12 1052 15
rect 1054 24 1062 26
rect 1054 22 1057 24
rect 1059 22 1062 24
rect 1054 12 1062 22
rect 1064 19 1069 26
rect 1096 20 1103 26
rect 1105 24 1113 26
rect 1105 22 1108 24
rect 1110 22 1113 24
rect 1105 20 1113 22
rect 1115 20 1123 26
rect 1064 16 1072 19
rect 1064 14 1067 16
rect 1069 14 1072 16
rect 1064 12 1072 14
rect 1067 9 1072 12
rect 1074 13 1082 19
rect 1074 11 1077 13
rect 1079 11 1082 13
rect 1074 9 1082 11
rect 1077 6 1082 9
rect 1084 17 1091 19
rect 1084 15 1087 17
rect 1089 15 1091 17
rect 1084 13 1091 15
rect 1096 13 1101 20
rect 1117 17 1123 20
rect 1125 24 1132 26
rect 1125 22 1128 24
rect 1130 22 1132 24
rect 1125 20 1132 22
rect 1125 17 1130 20
rect 1117 13 1121 17
rect 1084 6 1089 13
rect 1096 11 1102 13
rect 1096 9 1098 11
rect 1100 9 1102 11
rect 1096 7 1102 9
rect 1115 11 1121 13
rect 1115 9 1117 11
rect 1119 9 1121 11
rect 1115 7 1121 9
rect -145 -4 -136 -2
rect -145 -6 -142 -4
rect -140 -6 -136 -4
rect -145 -14 -136 -6
rect -93 -4 -84 -2
rect -93 -6 -90 -4
rect -88 -6 -84 -4
rect -93 -14 -84 -6
rect -41 -4 -32 -2
rect -41 -6 -38 -4
rect -36 -6 -32 -4
rect -41 -14 -32 -6
rect 11 -4 20 -2
rect 11 -6 14 -4
rect 16 -6 20 -4
rect 11 -14 20 -6
rect 63 -4 72 -2
rect 63 -6 66 -4
rect 68 -6 72 -4
rect 63 -14 72 -6
rect 116 -4 125 -2
rect 116 -6 119 -4
rect 121 -6 125 -4
rect 116 -14 125 -6
rect 304 -4 313 -2
rect 304 -6 307 -4
rect 309 -6 313 -4
rect 304 -14 313 -6
rect 357 -4 366 -2
rect 357 -6 360 -4
rect 362 -6 366 -4
rect 357 -14 366 -6
rect 409 -4 418 -2
rect 409 -6 412 -4
rect 414 -6 418 -4
rect 409 -14 418 -6
rect 461 -4 470 -2
rect 461 -6 464 -4
rect 466 -6 470 -4
rect 461 -14 470 -6
rect 513 -4 522 -2
rect 513 -6 516 -4
rect 518 -6 522 -4
rect 513 -14 522 -6
rect 612 -4 621 -2
rect 612 -6 615 -4
rect 617 -6 621 -4
rect 612 -14 621 -6
rect 665 -4 674 -2
rect 665 -6 668 -4
rect 670 -6 674 -4
rect 665 -14 674 -6
rect 717 -4 726 -2
rect 717 -6 720 -4
rect 722 -6 726 -4
rect 717 -14 726 -6
rect 769 -4 778 -2
rect 769 -6 772 -4
rect 774 -6 778 -4
rect 769 -14 778 -6
rect 821 -4 830 -2
rect 821 -6 824 -4
rect 826 -6 830 -4
rect 821 -14 830 -6
rect 873 -4 882 -2
rect 873 -6 876 -4
rect 878 -6 882 -4
rect 873 -14 882 -6
rect 926 -4 935 -2
rect 926 -6 929 -4
rect 931 -6 935 -4
rect 926 -14 935 -6
rect 980 -4 989 -2
rect 980 -6 983 -4
rect 985 -6 989 -4
rect 980 -14 989 -6
rect 1035 -4 1044 -2
rect 1035 -6 1038 -4
rect 1040 -6 1044 -4
rect 1035 -14 1044 -6
rect 1088 -4 1097 -2
rect 1088 -6 1091 -4
rect 1093 -6 1097 -4
rect 1088 -14 1097 -6
rect -145 -19 -134 -14
rect -156 -21 -149 -19
rect -156 -23 -154 -21
rect -152 -23 -149 -21
rect -156 -25 -149 -23
rect -147 -25 -134 -19
rect -132 -25 -127 -14
rect -125 -25 -120 -14
rect -118 -16 -111 -14
rect -118 -18 -115 -16
rect -113 -18 -111 -16
rect -118 -20 -111 -18
rect -93 -19 -82 -14
rect -118 -25 -113 -20
rect -104 -21 -97 -19
rect -104 -23 -102 -21
rect -100 -23 -97 -21
rect -104 -25 -97 -23
rect -95 -25 -82 -19
rect -80 -25 -75 -14
rect -73 -25 -68 -14
rect -66 -16 -59 -14
rect -66 -18 -63 -16
rect -61 -18 -59 -16
rect -66 -20 -59 -18
rect -41 -19 -30 -14
rect -66 -25 -61 -20
rect -52 -21 -45 -19
rect -52 -23 -50 -21
rect -48 -23 -45 -21
rect -52 -25 -45 -23
rect -43 -25 -30 -19
rect -28 -25 -23 -14
rect -21 -25 -16 -14
rect -14 -16 -7 -14
rect -14 -18 -11 -16
rect -9 -18 -7 -16
rect -14 -20 -7 -18
rect 11 -19 22 -14
rect -14 -25 -9 -20
rect 0 -21 7 -19
rect 0 -23 2 -21
rect 4 -23 7 -21
rect 0 -25 7 -23
rect 9 -25 22 -19
rect 24 -25 29 -14
rect 31 -25 36 -14
rect 38 -16 45 -14
rect 38 -18 41 -16
rect 43 -18 45 -16
rect 38 -20 45 -18
rect 63 -19 74 -14
rect 38 -25 43 -20
rect 52 -21 59 -19
rect 52 -23 54 -21
rect 56 -23 59 -21
rect 52 -25 59 -23
rect 61 -25 74 -19
rect 76 -25 81 -14
rect 83 -25 88 -14
rect 90 -16 97 -14
rect 90 -18 93 -16
rect 95 -18 97 -16
rect 90 -20 97 -18
rect 116 -19 127 -14
rect 90 -25 95 -20
rect 105 -21 112 -19
rect 105 -23 107 -21
rect 109 -23 112 -21
rect 105 -25 112 -23
rect 114 -25 127 -19
rect 129 -25 134 -14
rect 136 -25 141 -14
rect 143 -16 150 -14
rect 143 -18 146 -16
rect 148 -18 150 -16
rect 143 -20 150 -18
rect 304 -19 315 -14
rect 143 -25 148 -20
rect 162 -21 169 -19
rect 162 -23 164 -21
rect 166 -23 169 -21
rect 162 -25 169 -23
rect 171 -21 178 -19
rect 171 -23 174 -21
rect 176 -23 178 -21
rect 171 -25 178 -23
rect 182 -21 189 -19
rect 182 -23 184 -21
rect 186 -23 189 -21
rect 182 -25 189 -23
rect 191 -21 198 -19
rect 191 -23 194 -21
rect 196 -23 198 -21
rect 191 -25 198 -23
rect 202 -21 209 -19
rect 202 -23 204 -21
rect 206 -23 209 -21
rect 202 -25 209 -23
rect 211 -21 218 -19
rect 211 -23 214 -21
rect 216 -23 218 -21
rect 211 -25 218 -23
rect 224 -21 231 -19
rect 224 -23 226 -21
rect 228 -23 231 -21
rect 224 -25 231 -23
rect 233 -21 240 -19
rect 233 -23 236 -21
rect 238 -23 240 -21
rect 233 -25 240 -23
rect 246 -21 253 -19
rect 246 -23 248 -21
rect 250 -23 253 -21
rect 246 -25 253 -23
rect 255 -21 262 -19
rect 255 -23 258 -21
rect 260 -23 262 -21
rect 255 -25 262 -23
rect 268 -21 275 -19
rect 268 -23 270 -21
rect 272 -23 275 -21
rect 268 -25 275 -23
rect 277 -21 284 -19
rect 277 -23 280 -21
rect 282 -23 284 -21
rect 277 -25 284 -23
rect 293 -21 300 -19
rect 293 -23 295 -21
rect 297 -23 300 -21
rect 293 -25 300 -23
rect 302 -25 315 -19
rect 317 -25 322 -14
rect 324 -25 329 -14
rect 331 -16 338 -14
rect 331 -18 334 -16
rect 336 -18 338 -16
rect 331 -20 338 -18
rect 357 -19 368 -14
rect 331 -25 336 -20
rect 346 -21 353 -19
rect 346 -23 348 -21
rect 350 -23 353 -21
rect 346 -25 353 -23
rect 355 -25 368 -19
rect 370 -25 375 -14
rect 377 -25 382 -14
rect 384 -16 391 -14
rect 384 -18 387 -16
rect 389 -18 391 -16
rect 384 -20 391 -18
rect 409 -19 420 -14
rect 384 -25 389 -20
rect 398 -21 405 -19
rect 398 -23 400 -21
rect 402 -23 405 -21
rect 398 -25 405 -23
rect 407 -25 420 -19
rect 422 -25 427 -14
rect 429 -25 434 -14
rect 436 -16 443 -14
rect 436 -18 439 -16
rect 441 -18 443 -16
rect 436 -20 443 -18
rect 461 -19 472 -14
rect 436 -25 441 -20
rect 450 -21 457 -19
rect 450 -23 452 -21
rect 454 -23 457 -21
rect 450 -25 457 -23
rect 459 -25 472 -19
rect 474 -25 479 -14
rect 481 -25 486 -14
rect 488 -16 495 -14
rect 488 -18 491 -16
rect 493 -18 495 -16
rect 488 -20 495 -18
rect 513 -19 524 -14
rect 488 -25 493 -20
rect 502 -21 509 -19
rect 502 -23 504 -21
rect 506 -23 509 -21
rect 502 -25 509 -23
rect 511 -25 524 -19
rect 526 -25 531 -14
rect 533 -25 538 -14
rect 540 -16 547 -14
rect 540 -18 543 -16
rect 545 -18 547 -16
rect 540 -20 547 -18
rect 612 -19 623 -14
rect 540 -25 545 -20
rect 557 -21 564 -19
rect 557 -23 559 -21
rect 561 -23 564 -21
rect 557 -25 564 -23
rect 566 -21 573 -19
rect 566 -23 569 -21
rect 571 -23 573 -21
rect 566 -25 573 -23
rect 578 -21 585 -19
rect 578 -23 580 -21
rect 582 -23 585 -21
rect 578 -25 585 -23
rect 587 -21 594 -19
rect 587 -23 590 -21
rect 592 -23 594 -21
rect 587 -25 594 -23
rect 601 -21 608 -19
rect 601 -23 603 -21
rect 605 -23 608 -21
rect 601 -25 608 -23
rect 610 -25 623 -19
rect 625 -25 630 -14
rect 632 -25 637 -14
rect 639 -16 646 -14
rect 639 -18 642 -16
rect 644 -18 646 -16
rect 639 -20 646 -18
rect 665 -19 676 -14
rect 639 -25 644 -20
rect 654 -21 661 -19
rect 654 -23 656 -21
rect 658 -23 661 -21
rect 654 -25 661 -23
rect 663 -25 676 -19
rect 678 -25 683 -14
rect 685 -25 690 -14
rect 692 -16 699 -14
rect 692 -18 695 -16
rect 697 -18 699 -16
rect 692 -20 699 -18
rect 717 -19 728 -14
rect 692 -25 697 -20
rect 706 -21 713 -19
rect 706 -23 708 -21
rect 710 -23 713 -21
rect 706 -25 713 -23
rect 715 -25 728 -19
rect 730 -25 735 -14
rect 737 -25 742 -14
rect 744 -16 751 -14
rect 744 -18 747 -16
rect 749 -18 751 -16
rect 744 -20 751 -18
rect 769 -19 780 -14
rect 744 -25 749 -20
rect 758 -21 765 -19
rect 758 -23 760 -21
rect 762 -23 765 -21
rect 758 -25 765 -23
rect 767 -25 780 -19
rect 782 -25 787 -14
rect 789 -25 794 -14
rect 796 -16 803 -14
rect 796 -18 799 -16
rect 801 -18 803 -16
rect 796 -20 803 -18
rect 821 -19 832 -14
rect 796 -25 801 -20
rect 810 -21 817 -19
rect 810 -23 812 -21
rect 814 -23 817 -21
rect 810 -25 817 -23
rect 819 -25 832 -19
rect 834 -25 839 -14
rect 841 -25 846 -14
rect 848 -16 855 -14
rect 848 -18 851 -16
rect 853 -18 855 -16
rect 848 -20 855 -18
rect 873 -19 884 -14
rect 848 -25 853 -20
rect 862 -21 869 -19
rect 862 -23 864 -21
rect 866 -23 869 -21
rect 862 -25 869 -23
rect 871 -25 884 -19
rect 886 -25 891 -14
rect 893 -25 898 -14
rect 900 -16 907 -14
rect 900 -18 903 -16
rect 905 -18 907 -16
rect 900 -20 907 -18
rect 926 -19 937 -14
rect 900 -25 905 -20
rect 915 -21 922 -19
rect 915 -23 917 -21
rect 919 -23 922 -21
rect 915 -25 922 -23
rect 924 -25 937 -19
rect 939 -25 944 -14
rect 946 -25 951 -14
rect 953 -16 960 -14
rect 953 -18 956 -16
rect 958 -18 960 -16
rect 953 -20 960 -18
rect 980 -19 991 -14
rect 953 -25 958 -20
rect 969 -21 976 -19
rect 969 -23 971 -21
rect 973 -23 976 -21
rect 969 -25 976 -23
rect 978 -25 991 -19
rect 993 -25 998 -14
rect 1000 -25 1005 -14
rect 1007 -16 1014 -14
rect 1007 -18 1010 -16
rect 1012 -18 1014 -16
rect 1007 -20 1014 -18
rect 1035 -19 1046 -14
rect 1007 -25 1012 -20
rect 1024 -21 1031 -19
rect 1024 -23 1026 -21
rect 1028 -23 1031 -21
rect 1024 -25 1031 -23
rect 1033 -25 1046 -19
rect 1048 -25 1053 -14
rect 1055 -25 1060 -14
rect 1062 -16 1069 -14
rect 1062 -18 1065 -16
rect 1067 -18 1069 -16
rect 1062 -20 1069 -18
rect 1088 -19 1099 -14
rect 1062 -25 1067 -20
rect 1077 -21 1084 -19
rect 1077 -23 1079 -21
rect 1081 -23 1084 -21
rect 1077 -25 1084 -23
rect 1086 -25 1099 -19
rect 1101 -25 1106 -14
rect 1108 -25 1113 -14
rect 1115 -16 1122 -14
rect 1115 -18 1118 -16
rect 1120 -18 1122 -16
rect 1115 -20 1122 -18
rect 1115 -25 1120 -20
<< pdif >>
rect -273 333 -268 354
rect -275 331 -268 333
rect -275 329 -273 331
rect -271 329 -268 331
rect -275 327 -268 329
rect -266 352 -254 354
rect -266 350 -263 352
rect -261 350 -254 352
rect -266 345 -254 350
rect -237 345 -232 354
rect -266 343 -263 345
rect -261 343 -252 345
rect -266 327 -252 343
rect -250 338 -242 345
rect -250 336 -247 338
rect -245 336 -242 338
rect -250 331 -242 336
rect -250 329 -247 331
rect -245 329 -242 331
rect -250 327 -242 329
rect -240 338 -232 345
rect -240 336 -237 338
rect -235 336 -232 338
rect -240 327 -232 336
rect -230 348 -225 354
rect -230 346 -223 348
rect -230 344 -227 346
rect -225 344 -223 346
rect -230 342 -223 344
rect -213 342 -208 354
rect -230 327 -225 342
rect -215 340 -208 342
rect -215 338 -213 340
rect -211 338 -208 340
rect -215 333 -208 338
rect -215 331 -213 333
rect -211 331 -208 333
rect -215 329 -208 331
rect -206 352 -197 354
rect -206 350 -202 352
rect -200 350 -197 352
rect -174 352 -160 354
rect -174 351 -167 352
rect -206 342 -197 350
rect -190 342 -185 351
rect -206 329 -195 342
rect -193 333 -185 342
rect -193 331 -190 333
rect -188 331 -185 333
rect -193 329 -185 331
rect -190 326 -185 329
rect -183 326 -178 351
rect -176 350 -167 351
rect -165 350 -160 352
rect -176 345 -160 350
rect -176 343 -167 345
rect -165 343 -160 345
rect -176 326 -160 343
rect -158 344 -150 354
rect -158 342 -155 344
rect -153 342 -150 344
rect -158 337 -150 342
rect -158 335 -155 337
rect -153 335 -150 337
rect -158 326 -150 335
rect -148 352 -140 354
rect -148 350 -145 352
rect -143 350 -140 352
rect -148 345 -140 350
rect -148 343 -145 345
rect -143 343 -140 345
rect -148 326 -140 343
rect -138 339 -133 354
rect -123 339 -118 354
rect -138 337 -131 339
rect -138 335 -135 337
rect -133 335 -131 337
rect -138 330 -131 335
rect -138 328 -135 330
rect -133 328 -131 330
rect -138 326 -131 328
rect -125 337 -118 339
rect -125 335 -123 337
rect -121 335 -118 337
rect -125 330 -118 335
rect -125 328 -123 330
rect -121 328 -118 330
rect -125 326 -118 328
rect -116 352 -108 354
rect -116 350 -113 352
rect -111 350 -108 352
rect -116 345 -108 350
rect -116 343 -113 345
rect -111 343 -108 345
rect -116 326 -108 343
rect -106 344 -98 354
rect -106 342 -103 344
rect -101 342 -98 344
rect -106 337 -98 342
rect -106 335 -103 337
rect -101 335 -98 337
rect -106 326 -98 335
rect -96 352 -82 354
rect -96 350 -91 352
rect -89 351 -82 352
rect -59 352 -50 354
rect -89 350 -80 351
rect -96 345 -80 350
rect -96 343 -91 345
rect -89 343 -80 345
rect -96 326 -80 343
rect -78 326 -73 351
rect -71 342 -66 351
rect -59 350 -56 352
rect -54 350 -50 352
rect -59 342 -50 350
rect -71 333 -63 342
rect -71 331 -68 333
rect -66 331 -63 333
rect -71 329 -63 331
rect -61 329 -50 342
rect -48 342 -43 354
rect -34 347 -29 354
rect -36 345 -29 347
rect -36 343 -34 345
rect -32 343 -29 345
rect -48 340 -41 342
rect -36 341 -29 343
rect -48 338 -45 340
rect -43 338 -41 340
rect -48 333 -41 338
rect -34 333 -29 341
rect -27 333 -22 354
rect -20 352 -11 354
rect -20 350 -15 352
rect -13 350 -11 352
rect -20 344 -11 350
rect 7 345 14 347
rect -20 333 -9 344
rect -48 331 -45 333
rect -43 331 -41 333
rect -48 329 -41 331
rect -71 326 -66 329
rect -17 326 -9 333
rect -7 342 0 344
rect -7 340 -4 342
rect -2 340 0 342
rect -7 335 0 340
rect -7 333 -4 335
rect -2 333 0 335
rect 7 343 9 345
rect 11 343 14 345
rect 7 334 14 343
rect 16 345 24 347
rect 16 343 19 345
rect 21 343 24 345
rect 16 338 24 343
rect 16 336 19 338
rect 21 336 24 338
rect 16 334 24 336
rect 26 345 32 347
rect 47 345 54 347
rect 26 343 34 345
rect 26 341 29 343
rect 31 341 34 343
rect 26 334 34 341
rect -7 331 0 333
rect -7 326 -2 331
rect 28 327 34 334
rect 36 340 41 345
rect 47 343 49 345
rect 51 343 54 345
rect 36 338 43 340
rect 36 336 39 338
rect 41 336 43 338
rect 36 331 43 336
rect 47 334 54 343
rect 56 345 64 347
rect 56 343 59 345
rect 61 343 64 345
rect 56 338 64 343
rect 56 336 59 338
rect 61 336 64 338
rect 56 334 64 336
rect 66 345 72 347
rect 66 343 74 345
rect 66 341 69 343
rect 71 341 74 343
rect 66 334 74 341
rect 36 329 39 331
rect 41 329 43 331
rect 36 327 43 329
rect 68 327 74 334
rect 76 340 81 345
rect 89 342 94 354
rect 87 340 94 342
rect 76 338 83 340
rect 76 336 79 338
rect 81 336 83 338
rect 76 331 83 336
rect 76 329 79 331
rect 81 329 83 331
rect 87 338 89 340
rect 91 338 94 340
rect 87 333 94 338
rect 87 331 89 333
rect 91 331 94 333
rect 87 329 94 331
rect 96 352 105 354
rect 96 350 100 352
rect 102 350 105 352
rect 128 352 142 354
rect 128 351 135 352
rect 96 342 105 350
rect 112 342 117 351
rect 96 329 107 342
rect 109 333 117 342
rect 109 331 112 333
rect 114 331 117 333
rect 109 329 117 331
rect 76 327 83 329
rect 112 326 117 329
rect 119 326 124 351
rect 126 350 135 351
rect 137 350 142 352
rect 126 345 142 350
rect 126 343 135 345
rect 137 343 142 345
rect 126 326 142 343
rect 144 344 152 354
rect 144 342 147 344
rect 149 342 152 344
rect 144 337 152 342
rect 144 335 147 337
rect 149 335 152 337
rect 144 326 152 335
rect 154 352 162 354
rect 154 350 157 352
rect 159 350 162 352
rect 154 345 162 350
rect 154 343 157 345
rect 159 343 162 345
rect 154 326 162 343
rect 164 339 169 354
rect 179 339 184 354
rect 164 337 171 339
rect 164 335 167 337
rect 169 335 171 337
rect 164 330 171 335
rect 164 328 167 330
rect 169 328 171 330
rect 164 326 171 328
rect 177 337 184 339
rect 177 335 179 337
rect 181 335 184 337
rect 177 330 184 335
rect 177 328 179 330
rect 181 328 184 330
rect 177 326 184 328
rect 186 352 194 354
rect 186 350 189 352
rect 191 350 194 352
rect 186 345 194 350
rect 186 343 189 345
rect 191 343 194 345
rect 186 326 194 343
rect 196 344 204 354
rect 196 342 199 344
rect 201 342 204 344
rect 196 337 204 342
rect 196 335 199 337
rect 201 335 204 337
rect 196 326 204 335
rect 206 352 220 354
rect 206 350 211 352
rect 213 351 220 352
rect 243 352 252 354
rect 213 350 222 351
rect 206 345 222 350
rect 206 343 211 345
rect 213 343 222 345
rect 206 326 222 343
rect 224 326 229 351
rect 231 342 236 351
rect 243 350 246 352
rect 248 350 252 352
rect 243 342 252 350
rect 231 333 239 342
rect 231 331 234 333
rect 236 331 239 333
rect 231 329 239 331
rect 241 329 252 342
rect 254 342 259 354
rect 268 347 273 354
rect 266 345 273 347
rect 266 343 268 345
rect 270 343 273 345
rect 254 340 261 342
rect 266 341 273 343
rect 254 338 257 340
rect 259 338 261 340
rect 254 333 261 338
rect 268 333 273 341
rect 275 333 280 354
rect 282 352 291 354
rect 282 350 287 352
rect 289 350 291 352
rect 282 344 291 350
rect 314 345 321 347
rect 282 333 293 344
rect 254 331 257 333
rect 259 331 261 333
rect 254 329 261 331
rect 231 326 236 329
rect 285 326 293 333
rect 295 342 302 344
rect 295 340 298 342
rect 300 340 302 342
rect 295 335 302 340
rect 295 333 298 335
rect 300 333 302 335
rect 314 343 316 345
rect 318 343 321 345
rect 314 334 321 343
rect 323 345 331 347
rect 323 343 326 345
rect 328 343 331 345
rect 323 338 331 343
rect 323 336 326 338
rect 328 336 331 338
rect 323 334 331 336
rect 333 345 339 347
rect 333 343 341 345
rect 333 341 336 343
rect 338 341 341 343
rect 333 334 341 341
rect 295 331 302 333
rect 295 326 300 331
rect 335 327 341 334
rect 343 340 348 345
rect 366 342 371 354
rect 364 340 371 342
rect 343 338 350 340
rect 343 336 346 338
rect 348 336 350 338
rect 343 331 350 336
rect 343 329 346 331
rect 348 329 350 331
rect 364 338 366 340
rect 368 338 371 340
rect 364 333 371 338
rect 364 331 366 333
rect 368 331 371 333
rect 364 329 371 331
rect 373 352 382 354
rect 373 350 377 352
rect 379 350 382 352
rect 405 352 419 354
rect 405 351 412 352
rect 373 342 382 350
rect 389 342 394 351
rect 373 329 384 342
rect 386 333 394 342
rect 386 331 389 333
rect 391 331 394 333
rect 386 329 394 331
rect 343 327 350 329
rect 389 326 394 329
rect 396 326 401 351
rect 403 350 412 351
rect 414 350 419 352
rect 403 345 419 350
rect 403 343 412 345
rect 414 343 419 345
rect 403 326 419 343
rect 421 344 429 354
rect 421 342 424 344
rect 426 342 429 344
rect 421 337 429 342
rect 421 335 424 337
rect 426 335 429 337
rect 421 326 429 335
rect 431 352 439 354
rect 431 350 434 352
rect 436 350 439 352
rect 431 345 439 350
rect 431 343 434 345
rect 436 343 439 345
rect 431 326 439 343
rect 441 339 446 354
rect 456 339 461 354
rect 441 337 448 339
rect 441 335 444 337
rect 446 335 448 337
rect 441 330 448 335
rect 441 328 444 330
rect 446 328 448 330
rect 441 326 448 328
rect 454 337 461 339
rect 454 335 456 337
rect 458 335 461 337
rect 454 330 461 335
rect 454 328 456 330
rect 458 328 461 330
rect 454 326 461 328
rect 463 352 471 354
rect 463 350 466 352
rect 468 350 471 352
rect 463 345 471 350
rect 463 343 466 345
rect 468 343 471 345
rect 463 326 471 343
rect 473 344 481 354
rect 473 342 476 344
rect 478 342 481 344
rect 473 337 481 342
rect 473 335 476 337
rect 478 335 481 337
rect 473 326 481 335
rect 483 352 497 354
rect 483 350 488 352
rect 490 351 497 352
rect 520 352 529 354
rect 490 350 499 351
rect 483 345 499 350
rect 483 343 488 345
rect 490 343 499 345
rect 483 326 499 343
rect 501 326 506 351
rect 508 342 513 351
rect 520 350 523 352
rect 525 350 529 352
rect 520 342 529 350
rect 508 333 516 342
rect 508 331 511 333
rect 513 331 516 333
rect 508 329 516 331
rect 518 329 529 342
rect 531 342 536 354
rect 545 347 550 354
rect 543 345 550 347
rect 543 343 545 345
rect 547 343 550 345
rect 531 340 538 342
rect 543 341 550 343
rect 531 338 534 340
rect 536 338 538 340
rect 531 333 538 338
rect 545 333 550 341
rect 552 333 557 354
rect 559 352 568 354
rect 559 350 564 352
rect 566 350 568 352
rect 559 344 568 350
rect 591 345 598 347
rect 559 333 570 344
rect 531 331 534 333
rect 536 331 538 333
rect 531 329 538 331
rect 508 326 513 329
rect 562 326 570 333
rect 572 342 579 344
rect 572 340 575 342
rect 577 340 579 342
rect 572 335 579 340
rect 572 333 575 335
rect 577 333 579 335
rect 591 343 593 345
rect 595 343 598 345
rect 591 334 598 343
rect 600 345 608 347
rect 600 343 603 345
rect 605 343 608 345
rect 600 338 608 343
rect 600 336 603 338
rect 605 336 608 338
rect 600 334 608 336
rect 610 345 616 347
rect 610 343 618 345
rect 610 341 613 343
rect 615 341 618 343
rect 610 334 618 341
rect 572 331 579 333
rect 572 326 577 331
rect 612 327 618 334
rect 620 340 625 345
rect 642 342 647 354
rect 640 340 647 342
rect 620 338 627 340
rect 620 336 623 338
rect 625 336 627 338
rect 620 331 627 336
rect 620 329 623 331
rect 625 329 627 331
rect 640 338 642 340
rect 644 338 647 340
rect 640 333 647 338
rect 640 331 642 333
rect 644 331 647 333
rect 640 329 647 331
rect 649 352 658 354
rect 649 350 653 352
rect 655 350 658 352
rect 681 352 695 354
rect 681 351 688 352
rect 649 342 658 350
rect 665 342 670 351
rect 649 329 660 342
rect 662 333 670 342
rect 662 331 665 333
rect 667 331 670 333
rect 662 329 670 331
rect 620 327 627 329
rect 665 326 670 329
rect 672 326 677 351
rect 679 350 688 351
rect 690 350 695 352
rect 679 345 695 350
rect 679 343 688 345
rect 690 343 695 345
rect 679 326 695 343
rect 697 344 705 354
rect 697 342 700 344
rect 702 342 705 344
rect 697 337 705 342
rect 697 335 700 337
rect 702 335 705 337
rect 697 326 705 335
rect 707 352 715 354
rect 707 350 710 352
rect 712 350 715 352
rect 707 345 715 350
rect 707 343 710 345
rect 712 343 715 345
rect 707 326 715 343
rect 717 339 722 354
rect 732 339 737 354
rect 717 337 724 339
rect 717 335 720 337
rect 722 335 724 337
rect 717 330 724 335
rect 717 328 720 330
rect 722 328 724 330
rect 717 326 724 328
rect 730 337 737 339
rect 730 335 732 337
rect 734 335 737 337
rect 730 330 737 335
rect 730 328 732 330
rect 734 328 737 330
rect 730 326 737 328
rect 739 352 747 354
rect 739 350 742 352
rect 744 350 747 352
rect 739 345 747 350
rect 739 343 742 345
rect 744 343 747 345
rect 739 326 747 343
rect 749 344 757 354
rect 749 342 752 344
rect 754 342 757 344
rect 749 337 757 342
rect 749 335 752 337
rect 754 335 757 337
rect 749 326 757 335
rect 759 352 773 354
rect 759 350 764 352
rect 766 351 773 352
rect 796 352 805 354
rect 766 350 775 351
rect 759 345 775 350
rect 759 343 764 345
rect 766 343 775 345
rect 759 326 775 343
rect 777 326 782 351
rect 784 342 789 351
rect 796 350 799 352
rect 801 350 805 352
rect 796 342 805 350
rect 784 333 792 342
rect 784 331 787 333
rect 789 331 792 333
rect 784 329 792 331
rect 794 329 805 342
rect 807 342 812 354
rect 821 347 826 354
rect 819 345 826 347
rect 819 343 821 345
rect 823 343 826 345
rect 807 340 814 342
rect 819 341 826 343
rect 807 338 810 340
rect 812 338 814 340
rect 807 333 814 338
rect 821 333 826 341
rect 828 333 833 354
rect 835 352 844 354
rect 835 350 840 352
rect 842 350 844 352
rect 835 344 844 350
rect 867 345 874 347
rect 835 333 846 344
rect 807 331 810 333
rect 812 331 814 333
rect 807 329 814 331
rect 784 326 789 329
rect 838 326 846 333
rect 848 342 855 344
rect 848 340 851 342
rect 853 340 855 342
rect 848 335 855 340
rect 848 333 851 335
rect 853 333 855 335
rect 867 343 869 345
rect 871 343 874 345
rect 867 334 874 343
rect 876 345 884 347
rect 876 343 879 345
rect 881 343 884 345
rect 876 338 884 343
rect 876 336 879 338
rect 881 336 884 338
rect 876 334 884 336
rect 886 345 892 347
rect 886 343 894 345
rect 886 341 889 343
rect 891 341 894 343
rect 886 334 894 341
rect 848 331 855 333
rect 848 326 853 331
rect 888 327 894 334
rect 896 340 901 345
rect 919 342 924 354
rect 917 340 924 342
rect 896 338 903 340
rect 896 336 899 338
rect 901 336 903 338
rect 896 331 903 336
rect 896 329 899 331
rect 901 329 903 331
rect 917 338 919 340
rect 921 338 924 340
rect 917 333 924 338
rect 917 331 919 333
rect 921 331 924 333
rect 917 329 924 331
rect 926 352 935 354
rect 926 350 930 352
rect 932 350 935 352
rect 958 352 972 354
rect 958 351 965 352
rect 926 342 935 350
rect 942 342 947 351
rect 926 329 937 342
rect 939 333 947 342
rect 939 331 942 333
rect 944 331 947 333
rect 939 329 947 331
rect 896 327 903 329
rect 942 326 947 329
rect 949 326 954 351
rect 956 350 965 351
rect 967 350 972 352
rect 956 345 972 350
rect 956 343 965 345
rect 967 343 972 345
rect 956 326 972 343
rect 974 344 982 354
rect 974 342 977 344
rect 979 342 982 344
rect 974 337 982 342
rect 974 335 977 337
rect 979 335 982 337
rect 974 326 982 335
rect 984 352 992 354
rect 984 350 987 352
rect 989 350 992 352
rect 984 345 992 350
rect 984 343 987 345
rect 989 343 992 345
rect 984 326 992 343
rect 994 339 999 354
rect 1009 339 1014 354
rect 994 337 1001 339
rect 994 335 997 337
rect 999 335 1001 337
rect 994 330 1001 335
rect 994 328 997 330
rect 999 328 1001 330
rect 994 326 1001 328
rect 1007 337 1014 339
rect 1007 335 1009 337
rect 1011 335 1014 337
rect 1007 330 1014 335
rect 1007 328 1009 330
rect 1011 328 1014 330
rect 1007 326 1014 328
rect 1016 352 1024 354
rect 1016 350 1019 352
rect 1021 350 1024 352
rect 1016 345 1024 350
rect 1016 343 1019 345
rect 1021 343 1024 345
rect 1016 326 1024 343
rect 1026 344 1034 354
rect 1026 342 1029 344
rect 1031 342 1034 344
rect 1026 337 1034 342
rect 1026 335 1029 337
rect 1031 335 1034 337
rect 1026 326 1034 335
rect 1036 352 1050 354
rect 1036 350 1041 352
rect 1043 351 1050 352
rect 1073 352 1082 354
rect 1043 350 1052 351
rect 1036 345 1052 350
rect 1036 343 1041 345
rect 1043 343 1052 345
rect 1036 326 1052 343
rect 1054 326 1059 351
rect 1061 342 1066 351
rect 1073 350 1076 352
rect 1078 350 1082 352
rect 1073 342 1082 350
rect 1061 333 1069 342
rect 1061 331 1064 333
rect 1066 331 1069 333
rect 1061 329 1069 331
rect 1071 329 1082 342
rect 1084 342 1089 354
rect 1098 347 1103 354
rect 1096 345 1103 347
rect 1096 343 1098 345
rect 1100 343 1103 345
rect 1084 340 1091 342
rect 1096 341 1103 343
rect 1084 338 1087 340
rect 1089 338 1091 340
rect 1084 333 1091 338
rect 1098 333 1103 341
rect 1105 333 1110 354
rect 1112 352 1121 354
rect 1112 350 1117 352
rect 1119 350 1121 352
rect 1112 344 1121 350
rect 1112 333 1123 344
rect 1084 331 1087 333
rect 1089 331 1091 333
rect 1084 329 1091 331
rect 1061 326 1066 329
rect 1115 326 1123 333
rect 1125 342 1132 344
rect 1125 340 1128 342
rect 1130 340 1132 342
rect 1125 335 1132 340
rect 1125 333 1128 335
rect 1130 333 1132 335
rect 1125 331 1132 333
rect 1125 326 1130 331
rect -275 247 -268 249
rect -275 245 -273 247
rect -271 245 -268 247
rect -275 243 -268 245
rect -273 222 -268 243
rect -266 233 -252 249
rect -266 231 -263 233
rect -261 231 -252 233
rect -250 247 -242 249
rect -250 245 -247 247
rect -245 245 -242 247
rect -250 240 -242 245
rect -250 238 -247 240
rect -245 238 -242 240
rect -250 231 -242 238
rect -240 240 -232 249
rect -240 238 -237 240
rect -235 238 -232 240
rect -240 231 -232 238
rect -266 226 -254 231
rect -266 224 -263 226
rect -261 224 -254 226
rect -266 222 -254 224
rect -237 222 -232 231
rect -230 234 -225 249
rect -190 247 -185 250
rect -215 245 -208 247
rect -215 243 -213 245
rect -211 243 -208 245
rect -215 238 -208 243
rect -215 236 -213 238
rect -211 236 -208 238
rect -215 234 -208 236
rect -230 232 -223 234
rect -230 230 -227 232
rect -225 230 -223 232
rect -230 228 -223 230
rect -230 222 -225 228
rect -213 222 -208 234
rect -206 234 -195 247
rect -193 245 -185 247
rect -193 243 -190 245
rect -188 243 -185 245
rect -193 234 -185 243
rect -206 226 -197 234
rect -206 224 -202 226
rect -200 224 -197 226
rect -190 225 -185 234
rect -183 225 -178 250
rect -176 233 -160 250
rect -176 231 -167 233
rect -165 231 -160 233
rect -176 226 -160 231
rect -176 225 -167 226
rect -206 222 -197 224
rect -174 224 -167 225
rect -165 224 -160 226
rect -174 222 -160 224
rect -158 241 -150 250
rect -158 239 -155 241
rect -153 239 -150 241
rect -158 234 -150 239
rect -158 232 -155 234
rect -153 232 -150 234
rect -158 222 -150 232
rect -148 233 -140 250
rect -148 231 -145 233
rect -143 231 -140 233
rect -148 226 -140 231
rect -148 224 -145 226
rect -143 224 -140 226
rect -148 222 -140 224
rect -138 248 -131 250
rect -138 246 -135 248
rect -133 246 -131 248
rect -138 241 -131 246
rect -138 239 -135 241
rect -133 239 -131 241
rect -138 237 -131 239
rect -125 248 -118 250
rect -125 246 -123 248
rect -121 246 -118 248
rect -125 241 -118 246
rect -125 239 -123 241
rect -121 239 -118 241
rect -125 237 -118 239
rect -138 222 -133 237
rect -123 222 -118 237
rect -116 233 -108 250
rect -116 231 -113 233
rect -111 231 -108 233
rect -116 226 -108 231
rect -116 224 -113 226
rect -111 224 -108 226
rect -116 222 -108 224
rect -106 241 -98 250
rect -106 239 -103 241
rect -101 239 -98 241
rect -106 234 -98 239
rect -106 232 -103 234
rect -101 232 -98 234
rect -106 222 -98 232
rect -96 233 -80 250
rect -96 231 -91 233
rect -89 231 -80 233
rect -96 226 -80 231
rect -96 224 -91 226
rect -89 225 -80 226
rect -78 225 -73 250
rect -71 247 -66 250
rect -71 245 -63 247
rect -71 243 -68 245
rect -66 243 -63 245
rect -71 234 -63 243
rect -61 234 -50 247
rect -71 225 -66 234
rect -59 226 -50 234
rect -89 224 -82 225
rect -96 222 -82 224
rect -59 224 -56 226
rect -54 224 -50 226
rect -59 222 -50 224
rect -48 245 -41 247
rect -48 243 -45 245
rect -43 243 -41 245
rect -17 243 -9 250
rect -48 238 -41 243
rect -48 236 -45 238
rect -43 236 -41 238
rect -48 234 -41 236
rect -34 235 -29 243
rect -48 222 -43 234
rect -36 233 -29 235
rect -36 231 -34 233
rect -32 231 -29 233
rect -36 229 -29 231
rect -34 222 -29 229
rect -27 222 -22 243
rect -20 232 -9 243
rect -7 245 -2 250
rect -7 243 0 245
rect -7 241 -4 243
rect -2 241 0 243
rect 28 242 34 249
rect -7 236 0 241
rect -7 234 -4 236
rect -2 234 0 236
rect -7 232 0 234
rect 7 233 14 242
rect -20 226 -11 232
rect 7 231 9 233
rect 11 231 14 233
rect 7 229 14 231
rect 16 240 24 242
rect 16 238 19 240
rect 21 238 24 240
rect 16 233 24 238
rect 16 231 19 233
rect 21 231 24 233
rect 16 229 24 231
rect 26 235 34 242
rect 26 233 29 235
rect 31 233 34 235
rect 26 231 34 233
rect 36 246 43 249
rect 36 244 39 246
rect 41 244 43 246
rect 36 238 43 244
rect 68 242 74 249
rect 36 236 39 238
rect 41 236 43 238
rect 36 234 43 236
rect 36 231 41 234
rect 47 233 54 242
rect 47 231 49 233
rect 51 231 54 233
rect 26 229 32 231
rect -20 224 -15 226
rect -13 224 -11 226
rect -20 222 -11 224
rect 47 229 54 231
rect 56 240 64 242
rect 56 238 59 240
rect 61 238 64 240
rect 56 233 64 238
rect 56 231 59 233
rect 61 231 64 233
rect 56 229 64 231
rect 66 235 74 242
rect 66 233 69 235
rect 71 233 74 235
rect 66 231 74 233
rect 76 247 83 249
rect 112 247 117 250
rect 76 245 79 247
rect 81 245 83 247
rect 76 240 83 245
rect 76 238 79 240
rect 81 238 83 240
rect 76 236 83 238
rect 87 245 94 247
rect 87 243 89 245
rect 91 243 94 245
rect 87 238 94 243
rect 87 236 89 238
rect 91 236 94 238
rect 76 231 81 236
rect 87 234 94 236
rect 66 229 72 231
rect 89 222 94 234
rect 96 234 107 247
rect 109 245 117 247
rect 109 243 112 245
rect 114 243 117 245
rect 109 234 117 243
rect 96 226 105 234
rect 96 224 100 226
rect 102 224 105 226
rect 112 225 117 234
rect 119 225 124 250
rect 126 233 142 250
rect 126 231 135 233
rect 137 231 142 233
rect 126 226 142 231
rect 126 225 135 226
rect 96 222 105 224
rect 128 224 135 225
rect 137 224 142 226
rect 128 222 142 224
rect 144 241 152 250
rect 144 239 147 241
rect 149 239 152 241
rect 144 234 152 239
rect 144 232 147 234
rect 149 232 152 234
rect 144 222 152 232
rect 154 233 162 250
rect 154 231 157 233
rect 159 231 162 233
rect 154 226 162 231
rect 154 224 157 226
rect 159 224 162 226
rect 154 222 162 224
rect 164 248 171 250
rect 164 246 167 248
rect 169 246 171 248
rect 164 241 171 246
rect 164 239 167 241
rect 169 239 171 241
rect 164 237 171 239
rect 177 248 184 250
rect 177 246 179 248
rect 181 246 184 248
rect 177 241 184 246
rect 177 239 179 241
rect 181 239 184 241
rect 177 237 184 239
rect 164 222 169 237
rect 179 222 184 237
rect 186 233 194 250
rect 186 231 189 233
rect 191 231 194 233
rect 186 226 194 231
rect 186 224 189 226
rect 191 224 194 226
rect 186 222 194 224
rect 196 241 204 250
rect 196 239 199 241
rect 201 239 204 241
rect 196 234 204 239
rect 196 232 199 234
rect 201 232 204 234
rect 196 222 204 232
rect 206 233 222 250
rect 206 231 211 233
rect 213 231 222 233
rect 206 226 222 231
rect 206 224 211 226
rect 213 225 222 226
rect 224 225 229 250
rect 231 247 236 250
rect 231 245 239 247
rect 231 243 234 245
rect 236 243 239 245
rect 231 234 239 243
rect 241 234 252 247
rect 231 225 236 234
rect 243 226 252 234
rect 213 224 220 225
rect 206 222 220 224
rect 243 224 246 226
rect 248 224 252 226
rect 243 222 252 224
rect 254 245 261 247
rect 254 243 257 245
rect 259 243 261 245
rect 285 243 293 250
rect 254 238 261 243
rect 254 236 257 238
rect 259 236 261 238
rect 254 234 261 236
rect 268 235 273 243
rect 254 222 259 234
rect 266 233 273 235
rect 266 231 268 233
rect 270 231 273 233
rect 266 229 273 231
rect 268 222 273 229
rect 275 222 280 243
rect 282 232 293 243
rect 295 245 300 250
rect 295 243 302 245
rect 295 241 298 243
rect 300 241 302 243
rect 335 242 341 249
rect 295 236 302 241
rect 295 234 298 236
rect 300 234 302 236
rect 295 232 302 234
rect 314 233 321 242
rect 282 226 291 232
rect 314 231 316 233
rect 318 231 321 233
rect 314 229 321 231
rect 323 240 331 242
rect 323 238 326 240
rect 328 238 331 240
rect 323 233 331 238
rect 323 231 326 233
rect 328 231 331 233
rect 323 229 331 231
rect 333 235 341 242
rect 333 233 336 235
rect 338 233 341 235
rect 333 231 341 233
rect 343 247 350 249
rect 389 247 394 250
rect 343 245 346 247
rect 348 245 350 247
rect 343 240 350 245
rect 343 238 346 240
rect 348 238 350 240
rect 343 236 350 238
rect 364 245 371 247
rect 364 243 366 245
rect 368 243 371 245
rect 364 238 371 243
rect 364 236 366 238
rect 368 236 371 238
rect 343 231 348 236
rect 364 234 371 236
rect 333 229 339 231
rect 282 224 287 226
rect 289 224 291 226
rect 282 222 291 224
rect 366 222 371 234
rect 373 234 384 247
rect 386 245 394 247
rect 386 243 389 245
rect 391 243 394 245
rect 386 234 394 243
rect 373 226 382 234
rect 373 224 377 226
rect 379 224 382 226
rect 389 225 394 234
rect 396 225 401 250
rect 403 233 419 250
rect 403 231 412 233
rect 414 231 419 233
rect 403 226 419 231
rect 403 225 412 226
rect 373 222 382 224
rect 405 224 412 225
rect 414 224 419 226
rect 405 222 419 224
rect 421 241 429 250
rect 421 239 424 241
rect 426 239 429 241
rect 421 234 429 239
rect 421 232 424 234
rect 426 232 429 234
rect 421 222 429 232
rect 431 233 439 250
rect 431 231 434 233
rect 436 231 439 233
rect 431 226 439 231
rect 431 224 434 226
rect 436 224 439 226
rect 431 222 439 224
rect 441 248 448 250
rect 441 246 444 248
rect 446 246 448 248
rect 441 241 448 246
rect 441 239 444 241
rect 446 239 448 241
rect 441 237 448 239
rect 454 248 461 250
rect 454 246 456 248
rect 458 246 461 248
rect 454 241 461 246
rect 454 239 456 241
rect 458 239 461 241
rect 454 237 461 239
rect 441 222 446 237
rect 456 222 461 237
rect 463 233 471 250
rect 463 231 466 233
rect 468 231 471 233
rect 463 226 471 231
rect 463 224 466 226
rect 468 224 471 226
rect 463 222 471 224
rect 473 241 481 250
rect 473 239 476 241
rect 478 239 481 241
rect 473 234 481 239
rect 473 232 476 234
rect 478 232 481 234
rect 473 222 481 232
rect 483 233 499 250
rect 483 231 488 233
rect 490 231 499 233
rect 483 226 499 231
rect 483 224 488 226
rect 490 225 499 226
rect 501 225 506 250
rect 508 247 513 250
rect 508 245 516 247
rect 508 243 511 245
rect 513 243 516 245
rect 508 234 516 243
rect 518 234 529 247
rect 508 225 513 234
rect 520 226 529 234
rect 490 224 497 225
rect 483 222 497 224
rect 520 224 523 226
rect 525 224 529 226
rect 520 222 529 224
rect 531 245 538 247
rect 531 243 534 245
rect 536 243 538 245
rect 562 243 570 250
rect 531 238 538 243
rect 531 236 534 238
rect 536 236 538 238
rect 531 234 538 236
rect 545 235 550 243
rect 531 222 536 234
rect 543 233 550 235
rect 543 231 545 233
rect 547 231 550 233
rect 543 229 550 231
rect 545 222 550 229
rect 552 222 557 243
rect 559 232 570 243
rect 572 245 577 250
rect 572 243 579 245
rect 572 241 575 243
rect 577 241 579 243
rect 612 242 618 249
rect 572 236 579 241
rect 572 234 575 236
rect 577 234 579 236
rect 572 232 579 234
rect 591 233 598 242
rect 559 226 568 232
rect 591 231 593 233
rect 595 231 598 233
rect 591 229 598 231
rect 600 240 608 242
rect 600 238 603 240
rect 605 238 608 240
rect 600 233 608 238
rect 600 231 603 233
rect 605 231 608 233
rect 600 229 608 231
rect 610 235 618 242
rect 610 233 613 235
rect 615 233 618 235
rect 610 231 618 233
rect 620 247 627 249
rect 665 247 670 250
rect 620 245 623 247
rect 625 245 627 247
rect 620 240 627 245
rect 620 238 623 240
rect 625 238 627 240
rect 620 236 627 238
rect 640 245 647 247
rect 640 243 642 245
rect 644 243 647 245
rect 640 238 647 243
rect 640 236 642 238
rect 644 236 647 238
rect 620 231 625 236
rect 640 234 647 236
rect 610 229 616 231
rect 559 224 564 226
rect 566 224 568 226
rect 559 222 568 224
rect 642 222 647 234
rect 649 234 660 247
rect 662 245 670 247
rect 662 243 665 245
rect 667 243 670 245
rect 662 234 670 243
rect 649 226 658 234
rect 649 224 653 226
rect 655 224 658 226
rect 665 225 670 234
rect 672 225 677 250
rect 679 233 695 250
rect 679 231 688 233
rect 690 231 695 233
rect 679 226 695 231
rect 679 225 688 226
rect 649 222 658 224
rect 681 224 688 225
rect 690 224 695 226
rect 681 222 695 224
rect 697 241 705 250
rect 697 239 700 241
rect 702 239 705 241
rect 697 234 705 239
rect 697 232 700 234
rect 702 232 705 234
rect 697 222 705 232
rect 707 233 715 250
rect 707 231 710 233
rect 712 231 715 233
rect 707 226 715 231
rect 707 224 710 226
rect 712 224 715 226
rect 707 222 715 224
rect 717 248 724 250
rect 717 246 720 248
rect 722 246 724 248
rect 717 241 724 246
rect 717 239 720 241
rect 722 239 724 241
rect 717 237 724 239
rect 730 248 737 250
rect 730 246 732 248
rect 734 246 737 248
rect 730 241 737 246
rect 730 239 732 241
rect 734 239 737 241
rect 730 237 737 239
rect 717 222 722 237
rect 732 222 737 237
rect 739 233 747 250
rect 739 231 742 233
rect 744 231 747 233
rect 739 226 747 231
rect 739 224 742 226
rect 744 224 747 226
rect 739 222 747 224
rect 749 241 757 250
rect 749 239 752 241
rect 754 239 757 241
rect 749 234 757 239
rect 749 232 752 234
rect 754 232 757 234
rect 749 222 757 232
rect 759 233 775 250
rect 759 231 764 233
rect 766 231 775 233
rect 759 226 775 231
rect 759 224 764 226
rect 766 225 775 226
rect 777 225 782 250
rect 784 247 789 250
rect 784 245 792 247
rect 784 243 787 245
rect 789 243 792 245
rect 784 234 792 243
rect 794 234 805 247
rect 784 225 789 234
rect 796 226 805 234
rect 766 224 773 225
rect 759 222 773 224
rect 796 224 799 226
rect 801 224 805 226
rect 796 222 805 224
rect 807 245 814 247
rect 807 243 810 245
rect 812 243 814 245
rect 838 243 846 250
rect 807 238 814 243
rect 807 236 810 238
rect 812 236 814 238
rect 807 234 814 236
rect 821 235 826 243
rect 807 222 812 234
rect 819 233 826 235
rect 819 231 821 233
rect 823 231 826 233
rect 819 229 826 231
rect 821 222 826 229
rect 828 222 833 243
rect 835 232 846 243
rect 848 245 853 250
rect 848 243 855 245
rect 848 241 851 243
rect 853 241 855 243
rect 888 242 894 249
rect 848 236 855 241
rect 848 234 851 236
rect 853 234 855 236
rect 848 232 855 234
rect 867 233 874 242
rect 835 226 844 232
rect 867 231 869 233
rect 871 231 874 233
rect 867 229 874 231
rect 876 240 884 242
rect 876 238 879 240
rect 881 238 884 240
rect 876 233 884 238
rect 876 231 879 233
rect 881 231 884 233
rect 876 229 884 231
rect 886 235 894 242
rect 886 233 889 235
rect 891 233 894 235
rect 886 231 894 233
rect 896 247 903 249
rect 942 247 947 250
rect 896 245 899 247
rect 901 245 903 247
rect 896 240 903 245
rect 896 238 899 240
rect 901 238 903 240
rect 896 236 903 238
rect 917 245 924 247
rect 917 243 919 245
rect 921 243 924 245
rect 917 238 924 243
rect 917 236 919 238
rect 921 236 924 238
rect 896 231 901 236
rect 917 234 924 236
rect 886 229 892 231
rect 835 224 840 226
rect 842 224 844 226
rect 835 222 844 224
rect 919 222 924 234
rect 926 234 937 247
rect 939 245 947 247
rect 939 243 942 245
rect 944 243 947 245
rect 939 234 947 243
rect 926 226 935 234
rect 926 224 930 226
rect 932 224 935 226
rect 942 225 947 234
rect 949 225 954 250
rect 956 233 972 250
rect 956 231 965 233
rect 967 231 972 233
rect 956 226 972 231
rect 956 225 965 226
rect 926 222 935 224
rect 958 224 965 225
rect 967 224 972 226
rect 958 222 972 224
rect 974 241 982 250
rect 974 239 977 241
rect 979 239 982 241
rect 974 234 982 239
rect 974 232 977 234
rect 979 232 982 234
rect 974 222 982 232
rect 984 233 992 250
rect 984 231 987 233
rect 989 231 992 233
rect 984 226 992 231
rect 984 224 987 226
rect 989 224 992 226
rect 984 222 992 224
rect 994 248 1001 250
rect 994 246 997 248
rect 999 246 1001 248
rect 994 241 1001 246
rect 994 239 997 241
rect 999 239 1001 241
rect 994 237 1001 239
rect 1007 248 1014 250
rect 1007 246 1009 248
rect 1011 246 1014 248
rect 1007 241 1014 246
rect 1007 239 1009 241
rect 1011 239 1014 241
rect 1007 237 1014 239
rect 994 222 999 237
rect 1009 222 1014 237
rect 1016 233 1024 250
rect 1016 231 1019 233
rect 1021 231 1024 233
rect 1016 226 1024 231
rect 1016 224 1019 226
rect 1021 224 1024 226
rect 1016 222 1024 224
rect 1026 241 1034 250
rect 1026 239 1029 241
rect 1031 239 1034 241
rect 1026 234 1034 239
rect 1026 232 1029 234
rect 1031 232 1034 234
rect 1026 222 1034 232
rect 1036 233 1052 250
rect 1036 231 1041 233
rect 1043 231 1052 233
rect 1036 226 1052 231
rect 1036 224 1041 226
rect 1043 225 1052 226
rect 1054 225 1059 250
rect 1061 247 1066 250
rect 1061 245 1069 247
rect 1061 243 1064 245
rect 1066 243 1069 245
rect 1061 234 1069 243
rect 1071 234 1082 247
rect 1061 225 1066 234
rect 1073 226 1082 234
rect 1043 224 1050 225
rect 1036 222 1050 224
rect 1073 224 1076 226
rect 1078 224 1082 226
rect 1073 222 1082 224
rect 1084 245 1091 247
rect 1084 243 1087 245
rect 1089 243 1091 245
rect 1115 243 1123 250
rect 1084 238 1091 243
rect 1084 236 1087 238
rect 1089 236 1091 238
rect 1084 234 1091 236
rect 1098 235 1103 243
rect 1084 222 1089 234
rect 1096 233 1103 235
rect 1096 231 1098 233
rect 1100 231 1103 233
rect 1096 229 1103 231
rect 1098 222 1103 229
rect 1105 222 1110 243
rect 1112 232 1123 243
rect 1125 245 1130 250
rect 1125 243 1132 245
rect 1125 241 1128 243
rect 1130 241 1132 243
rect 1125 236 1132 241
rect 1125 234 1128 236
rect 1130 234 1132 236
rect 1125 232 1132 234
rect 1112 226 1121 232
rect 1112 224 1117 226
rect 1119 224 1121 226
rect 1112 222 1121 224
rect -273 189 -268 210
rect -275 187 -268 189
rect -275 185 -273 187
rect -271 185 -268 187
rect -275 183 -268 185
rect -266 208 -254 210
rect -266 206 -263 208
rect -261 206 -254 208
rect -266 201 -254 206
rect -237 201 -232 210
rect -266 199 -263 201
rect -261 199 -252 201
rect -266 183 -252 199
rect -250 194 -242 201
rect -250 192 -247 194
rect -245 192 -242 194
rect -250 187 -242 192
rect -250 185 -247 187
rect -245 185 -242 187
rect -250 183 -242 185
rect -240 194 -232 201
rect -240 192 -237 194
rect -235 192 -232 194
rect -240 183 -232 192
rect -230 204 -225 210
rect -230 202 -223 204
rect -230 200 -227 202
rect -225 200 -223 202
rect -230 198 -223 200
rect -213 198 -208 210
rect -230 183 -225 198
rect -215 196 -208 198
rect -215 194 -213 196
rect -211 194 -208 196
rect -215 189 -208 194
rect -215 187 -213 189
rect -211 187 -208 189
rect -215 185 -208 187
rect -206 208 -197 210
rect -206 206 -202 208
rect -200 206 -197 208
rect -174 208 -160 210
rect -174 207 -167 208
rect -206 198 -197 206
rect -190 198 -185 207
rect -206 185 -195 198
rect -193 189 -185 198
rect -193 187 -190 189
rect -188 187 -185 189
rect -193 185 -185 187
rect -190 182 -185 185
rect -183 182 -178 207
rect -176 206 -167 207
rect -165 206 -160 208
rect -176 201 -160 206
rect -176 199 -167 201
rect -165 199 -160 201
rect -176 182 -160 199
rect -158 200 -150 210
rect -158 198 -155 200
rect -153 198 -150 200
rect -158 193 -150 198
rect -158 191 -155 193
rect -153 191 -150 193
rect -158 182 -150 191
rect -148 208 -140 210
rect -148 206 -145 208
rect -143 206 -140 208
rect -148 201 -140 206
rect -148 199 -145 201
rect -143 199 -140 201
rect -148 182 -140 199
rect -138 195 -133 210
rect -123 195 -118 210
rect -138 193 -131 195
rect -138 191 -135 193
rect -133 191 -131 193
rect -138 186 -131 191
rect -138 184 -135 186
rect -133 184 -131 186
rect -138 182 -131 184
rect -125 193 -118 195
rect -125 191 -123 193
rect -121 191 -118 193
rect -125 186 -118 191
rect -125 184 -123 186
rect -121 184 -118 186
rect -125 182 -118 184
rect -116 208 -108 210
rect -116 206 -113 208
rect -111 206 -108 208
rect -116 201 -108 206
rect -116 199 -113 201
rect -111 199 -108 201
rect -116 182 -108 199
rect -106 200 -98 210
rect -106 198 -103 200
rect -101 198 -98 200
rect -106 193 -98 198
rect -106 191 -103 193
rect -101 191 -98 193
rect -106 182 -98 191
rect -96 208 -82 210
rect -96 206 -91 208
rect -89 207 -82 208
rect -59 208 -50 210
rect -89 206 -80 207
rect -96 201 -80 206
rect -96 199 -91 201
rect -89 199 -80 201
rect -96 182 -80 199
rect -78 182 -73 207
rect -71 198 -66 207
rect -59 206 -56 208
rect -54 206 -50 208
rect -59 198 -50 206
rect -71 189 -63 198
rect -71 187 -68 189
rect -66 187 -63 189
rect -71 185 -63 187
rect -61 185 -50 198
rect -48 198 -43 210
rect -34 203 -29 210
rect -36 201 -29 203
rect -36 199 -34 201
rect -32 199 -29 201
rect -48 196 -41 198
rect -36 197 -29 199
rect -48 194 -45 196
rect -43 194 -41 196
rect -48 189 -41 194
rect -34 189 -29 197
rect -27 189 -22 210
rect -20 208 -11 210
rect -20 206 -15 208
rect -13 206 -11 208
rect -20 200 -11 206
rect 7 201 14 203
rect -20 189 -9 200
rect -48 187 -45 189
rect -43 187 -41 189
rect -48 185 -41 187
rect -71 182 -66 185
rect -17 182 -9 189
rect -7 198 0 200
rect -7 196 -4 198
rect -2 196 0 198
rect -7 191 0 196
rect -7 189 -4 191
rect -2 189 0 191
rect 7 199 9 201
rect 11 199 14 201
rect 7 190 14 199
rect 16 201 24 203
rect 16 199 19 201
rect 21 199 24 201
rect 16 194 24 199
rect 16 192 19 194
rect 21 192 24 194
rect 16 190 24 192
rect 26 201 32 203
rect 47 201 54 203
rect 26 199 34 201
rect 26 197 29 199
rect 31 197 34 199
rect 26 190 34 197
rect -7 187 0 189
rect -7 182 -2 187
rect 28 183 34 190
rect 36 199 41 201
rect 47 199 49 201
rect 51 199 54 201
rect 36 197 43 199
rect 36 195 39 197
rect 41 195 43 197
rect 36 189 43 195
rect 47 190 54 199
rect 56 201 64 203
rect 56 199 59 201
rect 61 199 64 201
rect 56 194 64 199
rect 56 192 59 194
rect 61 192 64 194
rect 56 190 64 192
rect 66 201 72 203
rect 66 199 74 201
rect 66 197 69 199
rect 71 197 74 199
rect 66 190 74 197
rect 36 187 39 189
rect 41 187 43 189
rect 36 183 43 187
rect 68 183 74 190
rect 76 196 81 201
rect 89 198 94 210
rect 87 196 94 198
rect 76 194 83 196
rect 76 192 79 194
rect 81 192 83 194
rect 76 187 83 192
rect 76 185 79 187
rect 81 185 83 187
rect 87 194 89 196
rect 91 194 94 196
rect 87 189 94 194
rect 87 187 89 189
rect 91 187 94 189
rect 87 185 94 187
rect 96 208 105 210
rect 96 206 100 208
rect 102 206 105 208
rect 128 208 142 210
rect 128 207 135 208
rect 96 198 105 206
rect 112 198 117 207
rect 96 185 107 198
rect 109 189 117 198
rect 109 187 112 189
rect 114 187 117 189
rect 109 185 117 187
rect 76 183 83 185
rect 112 182 117 185
rect 119 182 124 207
rect 126 206 135 207
rect 137 206 142 208
rect 126 201 142 206
rect 126 199 135 201
rect 137 199 142 201
rect 126 182 142 199
rect 144 200 152 210
rect 144 198 147 200
rect 149 198 152 200
rect 144 193 152 198
rect 144 191 147 193
rect 149 191 152 193
rect 144 182 152 191
rect 154 208 162 210
rect 154 206 157 208
rect 159 206 162 208
rect 154 201 162 206
rect 154 199 157 201
rect 159 199 162 201
rect 154 182 162 199
rect 164 195 169 210
rect 179 195 184 210
rect 164 193 171 195
rect 164 191 167 193
rect 169 191 171 193
rect 164 186 171 191
rect 164 184 167 186
rect 169 184 171 186
rect 164 182 171 184
rect 177 193 184 195
rect 177 191 179 193
rect 181 191 184 193
rect 177 186 184 191
rect 177 184 179 186
rect 181 184 184 186
rect 177 182 184 184
rect 186 208 194 210
rect 186 206 189 208
rect 191 206 194 208
rect 186 201 194 206
rect 186 199 189 201
rect 191 199 194 201
rect 186 182 194 199
rect 196 200 204 210
rect 196 198 199 200
rect 201 198 204 200
rect 196 193 204 198
rect 196 191 199 193
rect 201 191 204 193
rect 196 182 204 191
rect 206 208 220 210
rect 206 206 211 208
rect 213 207 220 208
rect 243 208 252 210
rect 213 206 222 207
rect 206 201 222 206
rect 206 199 211 201
rect 213 199 222 201
rect 206 182 222 199
rect 224 182 229 207
rect 231 198 236 207
rect 243 206 246 208
rect 248 206 252 208
rect 243 198 252 206
rect 231 189 239 198
rect 231 187 234 189
rect 236 187 239 189
rect 231 185 239 187
rect 241 185 252 198
rect 254 198 259 210
rect 268 203 273 210
rect 266 201 273 203
rect 266 199 268 201
rect 270 199 273 201
rect 254 196 261 198
rect 266 197 273 199
rect 254 194 257 196
rect 259 194 261 196
rect 254 189 261 194
rect 268 189 273 197
rect 275 189 280 210
rect 282 208 291 210
rect 282 206 287 208
rect 289 206 291 208
rect 282 200 291 206
rect 314 201 321 203
rect 282 189 293 200
rect 254 187 257 189
rect 259 187 261 189
rect 254 185 261 187
rect 231 182 236 185
rect 285 182 293 189
rect 295 198 302 200
rect 295 196 298 198
rect 300 196 302 198
rect 295 191 302 196
rect 295 189 298 191
rect 300 189 302 191
rect 314 199 316 201
rect 318 199 321 201
rect 314 190 321 199
rect 323 201 331 203
rect 323 199 326 201
rect 328 199 331 201
rect 323 194 331 199
rect 323 192 326 194
rect 328 192 331 194
rect 323 190 331 192
rect 333 201 339 203
rect 333 199 341 201
rect 333 197 336 199
rect 338 197 341 199
rect 333 190 341 197
rect 295 187 302 189
rect 295 182 300 187
rect 335 183 341 190
rect 343 196 348 201
rect 366 198 371 210
rect 364 196 371 198
rect 343 194 350 196
rect 343 192 346 194
rect 348 192 350 194
rect 343 187 350 192
rect 343 185 346 187
rect 348 185 350 187
rect 364 194 366 196
rect 368 194 371 196
rect 364 189 371 194
rect 364 187 366 189
rect 368 187 371 189
rect 364 185 371 187
rect 373 208 382 210
rect 373 206 377 208
rect 379 206 382 208
rect 405 208 419 210
rect 405 207 412 208
rect 373 198 382 206
rect 389 198 394 207
rect 373 185 384 198
rect 386 189 394 198
rect 386 187 389 189
rect 391 187 394 189
rect 386 185 394 187
rect 343 183 350 185
rect 389 182 394 185
rect 396 182 401 207
rect 403 206 412 207
rect 414 206 419 208
rect 403 201 419 206
rect 403 199 412 201
rect 414 199 419 201
rect 403 182 419 199
rect 421 200 429 210
rect 421 198 424 200
rect 426 198 429 200
rect 421 193 429 198
rect 421 191 424 193
rect 426 191 429 193
rect 421 182 429 191
rect 431 208 439 210
rect 431 206 434 208
rect 436 206 439 208
rect 431 201 439 206
rect 431 199 434 201
rect 436 199 439 201
rect 431 182 439 199
rect 441 195 446 210
rect 456 195 461 210
rect 441 193 448 195
rect 441 191 444 193
rect 446 191 448 193
rect 441 186 448 191
rect 441 184 444 186
rect 446 184 448 186
rect 441 182 448 184
rect 454 193 461 195
rect 454 191 456 193
rect 458 191 461 193
rect 454 186 461 191
rect 454 184 456 186
rect 458 184 461 186
rect 454 182 461 184
rect 463 208 471 210
rect 463 206 466 208
rect 468 206 471 208
rect 463 201 471 206
rect 463 199 466 201
rect 468 199 471 201
rect 463 182 471 199
rect 473 200 481 210
rect 473 198 476 200
rect 478 198 481 200
rect 473 193 481 198
rect 473 191 476 193
rect 478 191 481 193
rect 473 182 481 191
rect 483 208 497 210
rect 483 206 488 208
rect 490 207 497 208
rect 520 208 529 210
rect 490 206 499 207
rect 483 201 499 206
rect 483 199 488 201
rect 490 199 499 201
rect 483 182 499 199
rect 501 182 506 207
rect 508 198 513 207
rect 520 206 523 208
rect 525 206 529 208
rect 520 198 529 206
rect 508 189 516 198
rect 508 187 511 189
rect 513 187 516 189
rect 508 185 516 187
rect 518 185 529 198
rect 531 198 536 210
rect 545 203 550 210
rect 543 201 550 203
rect 543 199 545 201
rect 547 199 550 201
rect 531 196 538 198
rect 543 197 550 199
rect 531 194 534 196
rect 536 194 538 196
rect 531 189 538 194
rect 545 189 550 197
rect 552 189 557 210
rect 559 208 568 210
rect 559 206 564 208
rect 566 206 568 208
rect 559 200 568 206
rect 591 201 598 203
rect 559 189 570 200
rect 531 187 534 189
rect 536 187 538 189
rect 531 185 538 187
rect 508 182 513 185
rect 562 182 570 189
rect 572 198 579 200
rect 572 196 575 198
rect 577 196 579 198
rect 572 191 579 196
rect 572 189 575 191
rect 577 189 579 191
rect 591 199 593 201
rect 595 199 598 201
rect 591 190 598 199
rect 600 201 608 203
rect 600 199 603 201
rect 605 199 608 201
rect 600 194 608 199
rect 600 192 603 194
rect 605 192 608 194
rect 600 190 608 192
rect 610 201 616 203
rect 610 199 618 201
rect 610 197 613 199
rect 615 197 618 199
rect 610 190 618 197
rect 572 187 579 189
rect 572 182 577 187
rect 612 183 618 190
rect 620 196 625 201
rect 642 198 647 210
rect 640 196 647 198
rect 620 194 627 196
rect 620 192 623 194
rect 625 192 627 194
rect 620 187 627 192
rect 620 185 623 187
rect 625 185 627 187
rect 640 194 642 196
rect 644 194 647 196
rect 640 189 647 194
rect 640 187 642 189
rect 644 187 647 189
rect 640 185 647 187
rect 649 208 658 210
rect 649 206 653 208
rect 655 206 658 208
rect 681 208 695 210
rect 681 207 688 208
rect 649 198 658 206
rect 665 198 670 207
rect 649 185 660 198
rect 662 189 670 198
rect 662 187 665 189
rect 667 187 670 189
rect 662 185 670 187
rect 620 183 627 185
rect 665 182 670 185
rect 672 182 677 207
rect 679 206 688 207
rect 690 206 695 208
rect 679 201 695 206
rect 679 199 688 201
rect 690 199 695 201
rect 679 182 695 199
rect 697 200 705 210
rect 697 198 700 200
rect 702 198 705 200
rect 697 193 705 198
rect 697 191 700 193
rect 702 191 705 193
rect 697 182 705 191
rect 707 208 715 210
rect 707 206 710 208
rect 712 206 715 208
rect 707 201 715 206
rect 707 199 710 201
rect 712 199 715 201
rect 707 182 715 199
rect 717 195 722 210
rect 732 195 737 210
rect 717 193 724 195
rect 717 191 720 193
rect 722 191 724 193
rect 717 186 724 191
rect 717 184 720 186
rect 722 184 724 186
rect 717 182 724 184
rect 730 193 737 195
rect 730 191 732 193
rect 734 191 737 193
rect 730 186 737 191
rect 730 184 732 186
rect 734 184 737 186
rect 730 182 737 184
rect 739 208 747 210
rect 739 206 742 208
rect 744 206 747 208
rect 739 201 747 206
rect 739 199 742 201
rect 744 199 747 201
rect 739 182 747 199
rect 749 200 757 210
rect 749 198 752 200
rect 754 198 757 200
rect 749 193 757 198
rect 749 191 752 193
rect 754 191 757 193
rect 749 182 757 191
rect 759 208 773 210
rect 759 206 764 208
rect 766 207 773 208
rect 796 208 805 210
rect 766 206 775 207
rect 759 201 775 206
rect 759 199 764 201
rect 766 199 775 201
rect 759 182 775 199
rect 777 182 782 207
rect 784 198 789 207
rect 796 206 799 208
rect 801 206 805 208
rect 796 198 805 206
rect 784 189 792 198
rect 784 187 787 189
rect 789 187 792 189
rect 784 185 792 187
rect 794 185 805 198
rect 807 198 812 210
rect 821 203 826 210
rect 819 201 826 203
rect 819 199 821 201
rect 823 199 826 201
rect 807 196 814 198
rect 819 197 826 199
rect 807 194 810 196
rect 812 194 814 196
rect 807 189 814 194
rect 821 189 826 197
rect 828 189 833 210
rect 835 208 844 210
rect 835 206 840 208
rect 842 206 844 208
rect 835 200 844 206
rect 867 201 874 203
rect 835 189 846 200
rect 807 187 810 189
rect 812 187 814 189
rect 807 185 814 187
rect 784 182 789 185
rect 838 182 846 189
rect 848 198 855 200
rect 848 196 851 198
rect 853 196 855 198
rect 848 191 855 196
rect 848 189 851 191
rect 853 189 855 191
rect 867 199 869 201
rect 871 199 874 201
rect 867 190 874 199
rect 876 201 884 203
rect 876 199 879 201
rect 881 199 884 201
rect 876 194 884 199
rect 876 192 879 194
rect 881 192 884 194
rect 876 190 884 192
rect 886 201 892 203
rect 886 199 894 201
rect 886 197 889 199
rect 891 197 894 199
rect 886 190 894 197
rect 848 187 855 189
rect 848 182 853 187
rect 888 183 894 190
rect 896 196 901 201
rect 919 198 924 210
rect 917 196 924 198
rect 896 194 903 196
rect 896 192 899 194
rect 901 192 903 194
rect 896 187 903 192
rect 896 185 899 187
rect 901 185 903 187
rect 917 194 919 196
rect 921 194 924 196
rect 917 189 924 194
rect 917 187 919 189
rect 921 187 924 189
rect 917 185 924 187
rect 926 208 935 210
rect 926 206 930 208
rect 932 206 935 208
rect 958 208 972 210
rect 958 207 965 208
rect 926 198 935 206
rect 942 198 947 207
rect 926 185 937 198
rect 939 189 947 198
rect 939 187 942 189
rect 944 187 947 189
rect 939 185 947 187
rect 896 183 903 185
rect 942 182 947 185
rect 949 182 954 207
rect 956 206 965 207
rect 967 206 972 208
rect 956 201 972 206
rect 956 199 965 201
rect 967 199 972 201
rect 956 182 972 199
rect 974 200 982 210
rect 974 198 977 200
rect 979 198 982 200
rect 974 193 982 198
rect 974 191 977 193
rect 979 191 982 193
rect 974 182 982 191
rect 984 208 992 210
rect 984 206 987 208
rect 989 206 992 208
rect 984 201 992 206
rect 984 199 987 201
rect 989 199 992 201
rect 984 182 992 199
rect 994 195 999 210
rect 1009 195 1014 210
rect 994 193 1001 195
rect 994 191 997 193
rect 999 191 1001 193
rect 994 186 1001 191
rect 994 184 997 186
rect 999 184 1001 186
rect 994 182 1001 184
rect 1007 193 1014 195
rect 1007 191 1009 193
rect 1011 191 1014 193
rect 1007 186 1014 191
rect 1007 184 1009 186
rect 1011 184 1014 186
rect 1007 182 1014 184
rect 1016 208 1024 210
rect 1016 206 1019 208
rect 1021 206 1024 208
rect 1016 201 1024 206
rect 1016 199 1019 201
rect 1021 199 1024 201
rect 1016 182 1024 199
rect 1026 200 1034 210
rect 1026 198 1029 200
rect 1031 198 1034 200
rect 1026 193 1034 198
rect 1026 191 1029 193
rect 1031 191 1034 193
rect 1026 182 1034 191
rect 1036 208 1050 210
rect 1036 206 1041 208
rect 1043 207 1050 208
rect 1073 208 1082 210
rect 1043 206 1052 207
rect 1036 201 1052 206
rect 1036 199 1041 201
rect 1043 199 1052 201
rect 1036 182 1052 199
rect 1054 182 1059 207
rect 1061 198 1066 207
rect 1073 206 1076 208
rect 1078 206 1082 208
rect 1073 198 1082 206
rect 1061 189 1069 198
rect 1061 187 1064 189
rect 1066 187 1069 189
rect 1061 185 1069 187
rect 1071 185 1082 198
rect 1084 198 1089 210
rect 1098 203 1103 210
rect 1096 201 1103 203
rect 1096 199 1098 201
rect 1100 199 1103 201
rect 1084 196 1091 198
rect 1096 197 1103 199
rect 1084 194 1087 196
rect 1089 194 1091 196
rect 1084 189 1091 194
rect 1098 189 1103 197
rect 1105 189 1110 210
rect 1112 208 1121 210
rect 1112 206 1117 208
rect 1119 206 1121 208
rect 1112 200 1121 206
rect 1112 189 1123 200
rect 1084 187 1087 189
rect 1089 187 1091 189
rect 1084 185 1091 187
rect 1061 182 1066 185
rect 1115 182 1123 189
rect 1125 198 1132 200
rect 1125 196 1128 198
rect 1130 196 1132 198
rect 1125 191 1132 196
rect 1125 189 1128 191
rect 1130 189 1132 191
rect 1125 187 1132 189
rect 1125 182 1130 187
rect -275 103 -268 105
rect -275 101 -273 103
rect -271 101 -268 103
rect -275 99 -268 101
rect -273 78 -268 99
rect -266 89 -252 105
rect -266 87 -263 89
rect -261 87 -252 89
rect -250 103 -242 105
rect -250 101 -247 103
rect -245 101 -242 103
rect -250 96 -242 101
rect -250 94 -247 96
rect -245 94 -242 96
rect -250 87 -242 94
rect -240 96 -232 105
rect -240 94 -237 96
rect -235 94 -232 96
rect -240 87 -232 94
rect -266 82 -254 87
rect -266 80 -263 82
rect -261 80 -254 82
rect -266 78 -254 80
rect -237 78 -232 87
rect -230 90 -225 105
rect -190 103 -185 106
rect -215 101 -208 103
rect -215 99 -213 101
rect -211 99 -208 101
rect -215 94 -208 99
rect -215 92 -213 94
rect -211 92 -208 94
rect -215 90 -208 92
rect -230 88 -223 90
rect -230 86 -227 88
rect -225 86 -223 88
rect -230 84 -223 86
rect -230 78 -225 84
rect -213 78 -208 90
rect -206 90 -195 103
rect -193 101 -185 103
rect -193 99 -190 101
rect -188 99 -185 101
rect -193 90 -185 99
rect -206 82 -197 90
rect -206 80 -202 82
rect -200 80 -197 82
rect -190 81 -185 90
rect -183 81 -178 106
rect -176 89 -160 106
rect -176 87 -167 89
rect -165 87 -160 89
rect -176 82 -160 87
rect -176 81 -167 82
rect -206 78 -197 80
rect -174 80 -167 81
rect -165 80 -160 82
rect -174 78 -160 80
rect -158 97 -150 106
rect -158 95 -155 97
rect -153 95 -150 97
rect -158 90 -150 95
rect -158 88 -155 90
rect -153 88 -150 90
rect -158 78 -150 88
rect -148 89 -140 106
rect -148 87 -145 89
rect -143 87 -140 89
rect -148 82 -140 87
rect -148 80 -145 82
rect -143 80 -140 82
rect -148 78 -140 80
rect -138 104 -131 106
rect -138 102 -135 104
rect -133 102 -131 104
rect -138 97 -131 102
rect -138 95 -135 97
rect -133 95 -131 97
rect -138 93 -131 95
rect -125 104 -118 106
rect -125 102 -123 104
rect -121 102 -118 104
rect -125 97 -118 102
rect -125 95 -123 97
rect -121 95 -118 97
rect -125 93 -118 95
rect -138 78 -133 93
rect -123 78 -118 93
rect -116 89 -108 106
rect -116 87 -113 89
rect -111 87 -108 89
rect -116 82 -108 87
rect -116 80 -113 82
rect -111 80 -108 82
rect -116 78 -108 80
rect -106 97 -98 106
rect -106 95 -103 97
rect -101 95 -98 97
rect -106 90 -98 95
rect -106 88 -103 90
rect -101 88 -98 90
rect -106 78 -98 88
rect -96 89 -80 106
rect -96 87 -91 89
rect -89 87 -80 89
rect -96 82 -80 87
rect -96 80 -91 82
rect -89 81 -80 82
rect -78 81 -73 106
rect -71 103 -66 106
rect -71 101 -63 103
rect -71 99 -68 101
rect -66 99 -63 101
rect -71 90 -63 99
rect -61 90 -50 103
rect -71 81 -66 90
rect -59 82 -50 90
rect -89 80 -82 81
rect -96 78 -82 80
rect -59 80 -56 82
rect -54 80 -50 82
rect -59 78 -50 80
rect -48 101 -41 103
rect -48 99 -45 101
rect -43 99 -41 101
rect -17 99 -9 106
rect -48 94 -41 99
rect -48 92 -45 94
rect -43 92 -41 94
rect -48 90 -41 92
rect -34 91 -29 99
rect -48 78 -43 90
rect -36 89 -29 91
rect -36 87 -34 89
rect -32 87 -29 89
rect -36 85 -29 87
rect -34 78 -29 85
rect -27 78 -22 99
rect -20 88 -9 99
rect -7 101 -2 106
rect -7 99 0 101
rect -7 97 -4 99
rect -2 97 0 99
rect 28 98 34 105
rect -7 92 0 97
rect -7 90 -4 92
rect -2 90 0 92
rect -7 88 0 90
rect 7 89 14 98
rect -20 82 -11 88
rect 7 87 9 89
rect 11 87 14 89
rect 7 85 14 87
rect 16 96 24 98
rect 16 94 19 96
rect 21 94 24 96
rect 16 89 24 94
rect 16 87 19 89
rect 21 87 24 89
rect 16 85 24 87
rect 26 91 34 98
rect 26 89 29 91
rect 31 89 34 91
rect 26 87 34 89
rect 36 100 43 105
rect 36 98 39 100
rect 41 98 43 100
rect 68 98 74 105
rect 36 93 43 98
rect 36 91 39 93
rect 41 91 43 93
rect 36 89 43 91
rect 47 89 54 98
rect 36 87 41 89
rect 47 87 49 89
rect 51 87 54 89
rect 26 85 32 87
rect -20 80 -15 82
rect -13 80 -11 82
rect -20 78 -11 80
rect 47 85 54 87
rect 56 96 64 98
rect 56 94 59 96
rect 61 94 64 96
rect 56 89 64 94
rect 56 87 59 89
rect 61 87 64 89
rect 56 85 64 87
rect 66 91 74 98
rect 66 89 69 91
rect 71 89 74 91
rect 66 87 74 89
rect 76 103 83 105
rect 112 103 117 106
rect 76 101 79 103
rect 81 101 83 103
rect 76 96 83 101
rect 76 94 79 96
rect 81 94 83 96
rect 76 92 83 94
rect 87 101 94 103
rect 87 99 89 101
rect 91 99 94 101
rect 87 94 94 99
rect 87 92 89 94
rect 91 92 94 94
rect 76 87 81 92
rect 87 90 94 92
rect 66 85 72 87
rect 89 78 94 90
rect 96 90 107 103
rect 109 101 117 103
rect 109 99 112 101
rect 114 99 117 101
rect 109 90 117 99
rect 96 82 105 90
rect 96 80 100 82
rect 102 80 105 82
rect 112 81 117 90
rect 119 81 124 106
rect 126 89 142 106
rect 126 87 135 89
rect 137 87 142 89
rect 126 82 142 87
rect 126 81 135 82
rect 96 78 105 80
rect 128 80 135 81
rect 137 80 142 82
rect 128 78 142 80
rect 144 97 152 106
rect 144 95 147 97
rect 149 95 152 97
rect 144 90 152 95
rect 144 88 147 90
rect 149 88 152 90
rect 144 78 152 88
rect 154 89 162 106
rect 154 87 157 89
rect 159 87 162 89
rect 154 82 162 87
rect 154 80 157 82
rect 159 80 162 82
rect 154 78 162 80
rect 164 104 171 106
rect 164 102 167 104
rect 169 102 171 104
rect 164 97 171 102
rect 164 95 167 97
rect 169 95 171 97
rect 164 93 171 95
rect 177 104 184 106
rect 177 102 179 104
rect 181 102 184 104
rect 177 97 184 102
rect 177 95 179 97
rect 181 95 184 97
rect 177 93 184 95
rect 164 78 169 93
rect 179 78 184 93
rect 186 89 194 106
rect 186 87 189 89
rect 191 87 194 89
rect 186 82 194 87
rect 186 80 189 82
rect 191 80 194 82
rect 186 78 194 80
rect 196 97 204 106
rect 196 95 199 97
rect 201 95 204 97
rect 196 90 204 95
rect 196 88 199 90
rect 201 88 204 90
rect 196 78 204 88
rect 206 89 222 106
rect 206 87 211 89
rect 213 87 222 89
rect 206 82 222 87
rect 206 80 211 82
rect 213 81 222 82
rect 224 81 229 106
rect 231 103 236 106
rect 231 101 239 103
rect 231 99 234 101
rect 236 99 239 101
rect 231 90 239 99
rect 241 90 252 103
rect 231 81 236 90
rect 243 82 252 90
rect 213 80 220 81
rect 206 78 220 80
rect 243 80 246 82
rect 248 80 252 82
rect 243 78 252 80
rect 254 101 261 103
rect 254 99 257 101
rect 259 99 261 101
rect 285 99 293 106
rect 254 94 261 99
rect 254 92 257 94
rect 259 92 261 94
rect 254 90 261 92
rect 268 91 273 99
rect 254 78 259 90
rect 266 89 273 91
rect 266 87 268 89
rect 270 87 273 89
rect 266 85 273 87
rect 268 78 273 85
rect 275 78 280 99
rect 282 88 293 99
rect 295 101 300 106
rect 295 99 302 101
rect 295 97 298 99
rect 300 97 302 99
rect 335 98 341 105
rect 295 92 302 97
rect 295 90 298 92
rect 300 90 302 92
rect 295 88 302 90
rect 314 89 321 98
rect 282 82 291 88
rect 314 87 316 89
rect 318 87 321 89
rect 314 85 321 87
rect 323 96 331 98
rect 323 94 326 96
rect 328 94 331 96
rect 323 89 331 94
rect 323 87 326 89
rect 328 87 331 89
rect 323 85 331 87
rect 333 91 341 98
rect 333 89 336 91
rect 338 89 341 91
rect 333 87 341 89
rect 343 103 350 105
rect 389 103 394 106
rect 343 101 346 103
rect 348 101 350 103
rect 343 96 350 101
rect 343 94 346 96
rect 348 94 350 96
rect 343 92 350 94
rect 364 101 371 103
rect 364 99 366 101
rect 368 99 371 101
rect 364 94 371 99
rect 364 92 366 94
rect 368 92 371 94
rect 343 87 348 92
rect 364 90 371 92
rect 333 85 339 87
rect 282 80 287 82
rect 289 80 291 82
rect 282 78 291 80
rect 366 78 371 90
rect 373 90 384 103
rect 386 101 394 103
rect 386 99 389 101
rect 391 99 394 101
rect 386 90 394 99
rect 373 82 382 90
rect 373 80 377 82
rect 379 80 382 82
rect 389 81 394 90
rect 396 81 401 106
rect 403 89 419 106
rect 403 87 412 89
rect 414 87 419 89
rect 403 82 419 87
rect 403 81 412 82
rect 373 78 382 80
rect 405 80 412 81
rect 414 80 419 82
rect 405 78 419 80
rect 421 97 429 106
rect 421 95 424 97
rect 426 95 429 97
rect 421 90 429 95
rect 421 88 424 90
rect 426 88 429 90
rect 421 78 429 88
rect 431 89 439 106
rect 431 87 434 89
rect 436 87 439 89
rect 431 82 439 87
rect 431 80 434 82
rect 436 80 439 82
rect 431 78 439 80
rect 441 104 448 106
rect 441 102 444 104
rect 446 102 448 104
rect 441 97 448 102
rect 441 95 444 97
rect 446 95 448 97
rect 441 93 448 95
rect 454 104 461 106
rect 454 102 456 104
rect 458 102 461 104
rect 454 97 461 102
rect 454 95 456 97
rect 458 95 461 97
rect 454 93 461 95
rect 441 78 446 93
rect 456 78 461 93
rect 463 89 471 106
rect 463 87 466 89
rect 468 87 471 89
rect 463 82 471 87
rect 463 80 466 82
rect 468 80 471 82
rect 463 78 471 80
rect 473 97 481 106
rect 473 95 476 97
rect 478 95 481 97
rect 473 90 481 95
rect 473 88 476 90
rect 478 88 481 90
rect 473 78 481 88
rect 483 89 499 106
rect 483 87 488 89
rect 490 87 499 89
rect 483 82 499 87
rect 483 80 488 82
rect 490 81 499 82
rect 501 81 506 106
rect 508 103 513 106
rect 508 101 516 103
rect 508 99 511 101
rect 513 99 516 101
rect 508 90 516 99
rect 518 90 529 103
rect 508 81 513 90
rect 520 82 529 90
rect 490 80 497 81
rect 483 78 497 80
rect 520 80 523 82
rect 525 80 529 82
rect 520 78 529 80
rect 531 101 538 103
rect 531 99 534 101
rect 536 99 538 101
rect 562 99 570 106
rect 531 94 538 99
rect 531 92 534 94
rect 536 92 538 94
rect 531 90 538 92
rect 545 91 550 99
rect 531 78 536 90
rect 543 89 550 91
rect 543 87 545 89
rect 547 87 550 89
rect 543 85 550 87
rect 545 78 550 85
rect 552 78 557 99
rect 559 88 570 99
rect 572 101 577 106
rect 572 99 579 101
rect 572 97 575 99
rect 577 97 579 99
rect 612 98 618 105
rect 572 92 579 97
rect 572 90 575 92
rect 577 90 579 92
rect 572 88 579 90
rect 591 89 598 98
rect 559 82 568 88
rect 591 87 593 89
rect 595 87 598 89
rect 591 85 598 87
rect 600 96 608 98
rect 600 94 603 96
rect 605 94 608 96
rect 600 89 608 94
rect 600 87 603 89
rect 605 87 608 89
rect 600 85 608 87
rect 610 91 618 98
rect 610 89 613 91
rect 615 89 618 91
rect 610 87 618 89
rect 620 103 627 105
rect 665 103 670 106
rect 620 101 623 103
rect 625 101 627 103
rect 620 96 627 101
rect 620 94 623 96
rect 625 94 627 96
rect 620 92 627 94
rect 640 101 647 103
rect 640 99 642 101
rect 644 99 647 101
rect 640 94 647 99
rect 640 92 642 94
rect 644 92 647 94
rect 620 87 625 92
rect 640 90 647 92
rect 610 85 616 87
rect 559 80 564 82
rect 566 80 568 82
rect 559 78 568 80
rect 642 78 647 90
rect 649 90 660 103
rect 662 101 670 103
rect 662 99 665 101
rect 667 99 670 101
rect 662 90 670 99
rect 649 82 658 90
rect 649 80 653 82
rect 655 80 658 82
rect 665 81 670 90
rect 672 81 677 106
rect 679 89 695 106
rect 679 87 688 89
rect 690 87 695 89
rect 679 82 695 87
rect 679 81 688 82
rect 649 78 658 80
rect 681 80 688 81
rect 690 80 695 82
rect 681 78 695 80
rect 697 97 705 106
rect 697 95 700 97
rect 702 95 705 97
rect 697 90 705 95
rect 697 88 700 90
rect 702 88 705 90
rect 697 78 705 88
rect 707 89 715 106
rect 707 87 710 89
rect 712 87 715 89
rect 707 82 715 87
rect 707 80 710 82
rect 712 80 715 82
rect 707 78 715 80
rect 717 104 724 106
rect 717 102 720 104
rect 722 102 724 104
rect 717 97 724 102
rect 717 95 720 97
rect 722 95 724 97
rect 717 93 724 95
rect 730 104 737 106
rect 730 102 732 104
rect 734 102 737 104
rect 730 97 737 102
rect 730 95 732 97
rect 734 95 737 97
rect 730 93 737 95
rect 717 78 722 93
rect 732 78 737 93
rect 739 89 747 106
rect 739 87 742 89
rect 744 87 747 89
rect 739 82 747 87
rect 739 80 742 82
rect 744 80 747 82
rect 739 78 747 80
rect 749 97 757 106
rect 749 95 752 97
rect 754 95 757 97
rect 749 90 757 95
rect 749 88 752 90
rect 754 88 757 90
rect 749 78 757 88
rect 759 89 775 106
rect 759 87 764 89
rect 766 87 775 89
rect 759 82 775 87
rect 759 80 764 82
rect 766 81 775 82
rect 777 81 782 106
rect 784 103 789 106
rect 784 101 792 103
rect 784 99 787 101
rect 789 99 792 101
rect 784 90 792 99
rect 794 90 805 103
rect 784 81 789 90
rect 796 82 805 90
rect 766 80 773 81
rect 759 78 773 80
rect 796 80 799 82
rect 801 80 805 82
rect 796 78 805 80
rect 807 101 814 103
rect 807 99 810 101
rect 812 99 814 101
rect 838 99 846 106
rect 807 94 814 99
rect 807 92 810 94
rect 812 92 814 94
rect 807 90 814 92
rect 821 91 826 99
rect 807 78 812 90
rect 819 89 826 91
rect 819 87 821 89
rect 823 87 826 89
rect 819 85 826 87
rect 821 78 826 85
rect 828 78 833 99
rect 835 88 846 99
rect 848 101 853 106
rect 848 99 855 101
rect 848 97 851 99
rect 853 97 855 99
rect 888 98 894 105
rect 848 92 855 97
rect 848 90 851 92
rect 853 90 855 92
rect 848 88 855 90
rect 867 89 874 98
rect 835 82 844 88
rect 867 87 869 89
rect 871 87 874 89
rect 867 85 874 87
rect 876 96 884 98
rect 876 94 879 96
rect 881 94 884 96
rect 876 89 884 94
rect 876 87 879 89
rect 881 87 884 89
rect 876 85 884 87
rect 886 91 894 98
rect 886 89 889 91
rect 891 89 894 91
rect 886 87 894 89
rect 896 103 903 105
rect 942 103 947 106
rect 896 101 899 103
rect 901 101 903 103
rect 896 96 903 101
rect 896 94 899 96
rect 901 94 903 96
rect 896 92 903 94
rect 917 101 924 103
rect 917 99 919 101
rect 921 99 924 101
rect 917 94 924 99
rect 917 92 919 94
rect 921 92 924 94
rect 896 87 901 92
rect 917 90 924 92
rect 886 85 892 87
rect 835 80 840 82
rect 842 80 844 82
rect 835 78 844 80
rect 919 78 924 90
rect 926 90 937 103
rect 939 101 947 103
rect 939 99 942 101
rect 944 99 947 101
rect 939 90 947 99
rect 926 82 935 90
rect 926 80 930 82
rect 932 80 935 82
rect 942 81 947 90
rect 949 81 954 106
rect 956 89 972 106
rect 956 87 965 89
rect 967 87 972 89
rect 956 82 972 87
rect 956 81 965 82
rect 926 78 935 80
rect 958 80 965 81
rect 967 80 972 82
rect 958 78 972 80
rect 974 97 982 106
rect 974 95 977 97
rect 979 95 982 97
rect 974 90 982 95
rect 974 88 977 90
rect 979 88 982 90
rect 974 78 982 88
rect 984 89 992 106
rect 984 87 987 89
rect 989 87 992 89
rect 984 82 992 87
rect 984 80 987 82
rect 989 80 992 82
rect 984 78 992 80
rect 994 104 1001 106
rect 994 102 997 104
rect 999 102 1001 104
rect 994 97 1001 102
rect 994 95 997 97
rect 999 95 1001 97
rect 994 93 1001 95
rect 1007 104 1014 106
rect 1007 102 1009 104
rect 1011 102 1014 104
rect 1007 97 1014 102
rect 1007 95 1009 97
rect 1011 95 1014 97
rect 1007 93 1014 95
rect 994 78 999 93
rect 1009 78 1014 93
rect 1016 89 1024 106
rect 1016 87 1019 89
rect 1021 87 1024 89
rect 1016 82 1024 87
rect 1016 80 1019 82
rect 1021 80 1024 82
rect 1016 78 1024 80
rect 1026 97 1034 106
rect 1026 95 1029 97
rect 1031 95 1034 97
rect 1026 90 1034 95
rect 1026 88 1029 90
rect 1031 88 1034 90
rect 1026 78 1034 88
rect 1036 89 1052 106
rect 1036 87 1041 89
rect 1043 87 1052 89
rect 1036 82 1052 87
rect 1036 80 1041 82
rect 1043 81 1052 82
rect 1054 81 1059 106
rect 1061 103 1066 106
rect 1061 101 1069 103
rect 1061 99 1064 101
rect 1066 99 1069 101
rect 1061 90 1069 99
rect 1071 90 1082 103
rect 1061 81 1066 90
rect 1073 82 1082 90
rect 1043 80 1050 81
rect 1036 78 1050 80
rect 1073 80 1076 82
rect 1078 80 1082 82
rect 1073 78 1082 80
rect 1084 101 1091 103
rect 1084 99 1087 101
rect 1089 99 1091 101
rect 1115 99 1123 106
rect 1084 94 1091 99
rect 1084 92 1087 94
rect 1089 92 1091 94
rect 1084 90 1091 92
rect 1098 91 1103 99
rect 1084 78 1089 90
rect 1096 89 1103 91
rect 1096 87 1098 89
rect 1100 87 1103 89
rect 1096 85 1103 87
rect 1098 78 1103 85
rect 1105 78 1110 99
rect 1112 88 1123 99
rect 1125 101 1130 106
rect 1125 99 1132 101
rect 1125 97 1128 99
rect 1130 97 1132 99
rect 1125 92 1132 97
rect 1125 90 1128 92
rect 1130 90 1132 92
rect 1125 88 1132 90
rect 1112 82 1121 88
rect 1112 80 1117 82
rect 1119 80 1121 82
rect 1112 78 1121 80
rect -273 45 -268 66
rect -275 43 -268 45
rect -275 41 -273 43
rect -271 41 -268 43
rect -275 39 -268 41
rect -266 64 -254 66
rect -266 62 -263 64
rect -261 62 -254 64
rect -266 57 -254 62
rect -237 57 -232 66
rect -266 55 -263 57
rect -261 55 -252 57
rect -266 39 -252 55
rect -250 50 -242 57
rect -250 48 -247 50
rect -245 48 -242 50
rect -250 43 -242 48
rect -250 41 -247 43
rect -245 41 -242 43
rect -250 39 -242 41
rect -240 50 -232 57
rect -240 48 -237 50
rect -235 48 -232 50
rect -240 39 -232 48
rect -230 60 -225 66
rect -230 58 -223 60
rect -230 56 -227 58
rect -225 56 -223 58
rect -230 54 -223 56
rect -213 54 -208 66
rect -230 39 -225 54
rect -215 52 -208 54
rect -215 50 -213 52
rect -211 50 -208 52
rect -215 45 -208 50
rect -215 43 -213 45
rect -211 43 -208 45
rect -215 41 -208 43
rect -206 64 -197 66
rect -206 62 -202 64
rect -200 62 -197 64
rect -174 64 -160 66
rect -174 63 -167 64
rect -206 54 -197 62
rect -190 54 -185 63
rect -206 41 -195 54
rect -193 45 -185 54
rect -193 43 -190 45
rect -188 43 -185 45
rect -193 41 -185 43
rect -190 38 -185 41
rect -183 38 -178 63
rect -176 62 -167 63
rect -165 62 -160 64
rect -176 57 -160 62
rect -176 55 -167 57
rect -165 55 -160 57
rect -176 38 -160 55
rect -158 56 -150 66
rect -158 54 -155 56
rect -153 54 -150 56
rect -158 49 -150 54
rect -158 47 -155 49
rect -153 47 -150 49
rect -158 38 -150 47
rect -148 64 -140 66
rect -148 62 -145 64
rect -143 62 -140 64
rect -148 57 -140 62
rect -148 55 -145 57
rect -143 55 -140 57
rect -148 38 -140 55
rect -138 51 -133 66
rect -123 51 -118 66
rect -138 49 -131 51
rect -138 47 -135 49
rect -133 47 -131 49
rect -138 42 -131 47
rect -138 40 -135 42
rect -133 40 -131 42
rect -138 38 -131 40
rect -125 49 -118 51
rect -125 47 -123 49
rect -121 47 -118 49
rect -125 42 -118 47
rect -125 40 -123 42
rect -121 40 -118 42
rect -125 38 -118 40
rect -116 64 -108 66
rect -116 62 -113 64
rect -111 62 -108 64
rect -116 57 -108 62
rect -116 55 -113 57
rect -111 55 -108 57
rect -116 38 -108 55
rect -106 56 -98 66
rect -106 54 -103 56
rect -101 54 -98 56
rect -106 49 -98 54
rect -106 47 -103 49
rect -101 47 -98 49
rect -106 38 -98 47
rect -96 64 -82 66
rect -96 62 -91 64
rect -89 63 -82 64
rect -59 64 -50 66
rect -89 62 -80 63
rect -96 57 -80 62
rect -96 55 -91 57
rect -89 55 -80 57
rect -96 38 -80 55
rect -78 38 -73 63
rect -71 54 -66 63
rect -59 62 -56 64
rect -54 62 -50 64
rect -59 54 -50 62
rect -71 45 -63 54
rect -71 43 -68 45
rect -66 43 -63 45
rect -71 41 -63 43
rect -61 41 -50 54
rect -48 54 -43 66
rect -34 59 -29 66
rect -36 57 -29 59
rect -36 55 -34 57
rect -32 55 -29 57
rect -48 52 -41 54
rect -36 53 -29 55
rect -48 50 -45 52
rect -43 50 -41 52
rect -48 45 -41 50
rect -34 45 -29 53
rect -27 45 -22 66
rect -20 64 -11 66
rect -20 62 -15 64
rect -13 62 -11 64
rect -20 56 -11 62
rect 7 57 14 59
rect -20 45 -9 56
rect -48 43 -45 45
rect -43 43 -41 45
rect -48 41 -41 43
rect -71 38 -66 41
rect -17 38 -9 45
rect -7 54 0 56
rect -7 52 -4 54
rect -2 52 0 54
rect -7 47 0 52
rect -7 45 -4 47
rect -2 45 0 47
rect 7 55 9 57
rect 11 55 14 57
rect 7 46 14 55
rect 16 57 24 59
rect 16 55 19 57
rect 21 55 24 57
rect 16 50 24 55
rect 16 48 19 50
rect 21 48 24 50
rect 16 46 24 48
rect 26 57 32 59
rect 47 57 54 59
rect 26 55 34 57
rect 26 53 29 55
rect 31 53 34 55
rect 26 46 34 53
rect -7 43 0 45
rect -7 38 -2 43
rect 28 39 34 46
rect 36 52 41 57
rect 47 55 49 57
rect 51 55 54 57
rect 36 50 43 52
rect 36 48 39 50
rect 41 48 43 50
rect 36 43 43 48
rect 47 46 54 55
rect 56 57 64 59
rect 56 55 59 57
rect 61 55 64 57
rect 56 50 64 55
rect 56 48 59 50
rect 61 48 64 50
rect 56 46 64 48
rect 66 57 72 59
rect 66 55 74 57
rect 66 53 69 55
rect 71 53 74 55
rect 66 46 74 53
rect 36 41 39 43
rect 41 41 43 43
rect 36 39 43 41
rect 68 39 74 46
rect 76 52 81 57
rect 89 54 94 66
rect 87 52 94 54
rect 76 50 83 52
rect 76 48 79 50
rect 81 48 83 50
rect 76 43 83 48
rect 76 41 79 43
rect 81 41 83 43
rect 87 50 89 52
rect 91 50 94 52
rect 87 45 94 50
rect 87 43 89 45
rect 91 43 94 45
rect 87 41 94 43
rect 96 64 105 66
rect 96 62 100 64
rect 102 62 105 64
rect 128 64 142 66
rect 128 63 135 64
rect 96 54 105 62
rect 112 54 117 63
rect 96 41 107 54
rect 109 45 117 54
rect 109 43 112 45
rect 114 43 117 45
rect 109 41 117 43
rect 76 39 83 41
rect 112 38 117 41
rect 119 38 124 63
rect 126 62 135 63
rect 137 62 142 64
rect 126 57 142 62
rect 126 55 135 57
rect 137 55 142 57
rect 126 38 142 55
rect 144 56 152 66
rect 144 54 147 56
rect 149 54 152 56
rect 144 49 152 54
rect 144 47 147 49
rect 149 47 152 49
rect 144 38 152 47
rect 154 64 162 66
rect 154 62 157 64
rect 159 62 162 64
rect 154 57 162 62
rect 154 55 157 57
rect 159 55 162 57
rect 154 38 162 55
rect 164 51 169 66
rect 179 51 184 66
rect 164 49 171 51
rect 164 47 167 49
rect 169 47 171 49
rect 164 42 171 47
rect 164 40 167 42
rect 169 40 171 42
rect 164 38 171 40
rect 177 49 184 51
rect 177 47 179 49
rect 181 47 184 49
rect 177 42 184 47
rect 177 40 179 42
rect 181 40 184 42
rect 177 38 184 40
rect 186 64 194 66
rect 186 62 189 64
rect 191 62 194 64
rect 186 57 194 62
rect 186 55 189 57
rect 191 55 194 57
rect 186 38 194 55
rect 196 56 204 66
rect 196 54 199 56
rect 201 54 204 56
rect 196 49 204 54
rect 196 47 199 49
rect 201 47 204 49
rect 196 38 204 47
rect 206 64 220 66
rect 206 62 211 64
rect 213 63 220 64
rect 243 64 252 66
rect 213 62 222 63
rect 206 57 222 62
rect 206 55 211 57
rect 213 55 222 57
rect 206 38 222 55
rect 224 38 229 63
rect 231 54 236 63
rect 243 62 246 64
rect 248 62 252 64
rect 243 54 252 62
rect 231 45 239 54
rect 231 43 234 45
rect 236 43 239 45
rect 231 41 239 43
rect 241 41 252 54
rect 254 54 259 66
rect 268 59 273 66
rect 266 57 273 59
rect 266 55 268 57
rect 270 55 273 57
rect 254 52 261 54
rect 266 53 273 55
rect 254 50 257 52
rect 259 50 261 52
rect 254 45 261 50
rect 268 45 273 53
rect 275 45 280 66
rect 282 64 291 66
rect 282 62 287 64
rect 289 62 291 64
rect 282 56 291 62
rect 314 57 321 59
rect 282 45 293 56
rect 254 43 257 45
rect 259 43 261 45
rect 254 41 261 43
rect 231 38 236 41
rect 285 38 293 45
rect 295 54 302 56
rect 295 52 298 54
rect 300 52 302 54
rect 295 47 302 52
rect 295 45 298 47
rect 300 45 302 47
rect 314 55 316 57
rect 318 55 321 57
rect 314 46 321 55
rect 323 57 331 59
rect 323 55 326 57
rect 328 55 331 57
rect 323 50 331 55
rect 323 48 326 50
rect 328 48 331 50
rect 323 46 331 48
rect 333 57 339 59
rect 333 55 341 57
rect 333 53 336 55
rect 338 53 341 55
rect 333 46 341 53
rect 295 43 302 45
rect 295 38 300 43
rect 335 39 341 46
rect 343 52 348 57
rect 366 54 371 66
rect 364 52 371 54
rect 343 50 350 52
rect 343 48 346 50
rect 348 48 350 50
rect 343 43 350 48
rect 343 41 346 43
rect 348 41 350 43
rect 364 50 366 52
rect 368 50 371 52
rect 364 45 371 50
rect 364 43 366 45
rect 368 43 371 45
rect 364 41 371 43
rect 373 64 382 66
rect 373 62 377 64
rect 379 62 382 64
rect 405 64 419 66
rect 405 63 412 64
rect 373 54 382 62
rect 389 54 394 63
rect 373 41 384 54
rect 386 45 394 54
rect 386 43 389 45
rect 391 43 394 45
rect 386 41 394 43
rect 343 39 350 41
rect 389 38 394 41
rect 396 38 401 63
rect 403 62 412 63
rect 414 62 419 64
rect 403 57 419 62
rect 403 55 412 57
rect 414 55 419 57
rect 403 38 419 55
rect 421 56 429 66
rect 421 54 424 56
rect 426 54 429 56
rect 421 49 429 54
rect 421 47 424 49
rect 426 47 429 49
rect 421 38 429 47
rect 431 64 439 66
rect 431 62 434 64
rect 436 62 439 64
rect 431 57 439 62
rect 431 55 434 57
rect 436 55 439 57
rect 431 38 439 55
rect 441 51 446 66
rect 456 51 461 66
rect 441 49 448 51
rect 441 47 444 49
rect 446 47 448 49
rect 441 42 448 47
rect 441 40 444 42
rect 446 40 448 42
rect 441 38 448 40
rect 454 49 461 51
rect 454 47 456 49
rect 458 47 461 49
rect 454 42 461 47
rect 454 40 456 42
rect 458 40 461 42
rect 454 38 461 40
rect 463 64 471 66
rect 463 62 466 64
rect 468 62 471 64
rect 463 57 471 62
rect 463 55 466 57
rect 468 55 471 57
rect 463 38 471 55
rect 473 56 481 66
rect 473 54 476 56
rect 478 54 481 56
rect 473 49 481 54
rect 473 47 476 49
rect 478 47 481 49
rect 473 38 481 47
rect 483 64 497 66
rect 483 62 488 64
rect 490 63 497 64
rect 520 64 529 66
rect 490 62 499 63
rect 483 57 499 62
rect 483 55 488 57
rect 490 55 499 57
rect 483 38 499 55
rect 501 38 506 63
rect 508 54 513 63
rect 520 62 523 64
rect 525 62 529 64
rect 520 54 529 62
rect 508 45 516 54
rect 508 43 511 45
rect 513 43 516 45
rect 508 41 516 43
rect 518 41 529 54
rect 531 54 536 66
rect 545 59 550 66
rect 543 57 550 59
rect 543 55 545 57
rect 547 55 550 57
rect 531 52 538 54
rect 543 53 550 55
rect 531 50 534 52
rect 536 50 538 52
rect 531 45 538 50
rect 545 45 550 53
rect 552 45 557 66
rect 559 64 568 66
rect 559 62 564 64
rect 566 62 568 64
rect 559 56 568 62
rect 591 57 598 59
rect 559 45 570 56
rect 531 43 534 45
rect 536 43 538 45
rect 531 41 538 43
rect 508 38 513 41
rect 562 38 570 45
rect 572 54 579 56
rect 572 52 575 54
rect 577 52 579 54
rect 572 47 579 52
rect 572 45 575 47
rect 577 45 579 47
rect 591 55 593 57
rect 595 55 598 57
rect 591 46 598 55
rect 600 57 608 59
rect 600 55 603 57
rect 605 55 608 57
rect 600 50 608 55
rect 600 48 603 50
rect 605 48 608 50
rect 600 46 608 48
rect 610 57 616 59
rect 610 55 618 57
rect 610 53 613 55
rect 615 53 618 55
rect 610 46 618 53
rect 572 43 579 45
rect 572 38 577 43
rect 612 39 618 46
rect 620 52 625 57
rect 642 54 647 66
rect 640 52 647 54
rect 620 50 627 52
rect 620 48 623 50
rect 625 48 627 50
rect 620 43 627 48
rect 620 41 623 43
rect 625 41 627 43
rect 640 50 642 52
rect 644 50 647 52
rect 640 45 647 50
rect 640 43 642 45
rect 644 43 647 45
rect 640 41 647 43
rect 649 64 658 66
rect 649 62 653 64
rect 655 62 658 64
rect 681 64 695 66
rect 681 63 688 64
rect 649 54 658 62
rect 665 54 670 63
rect 649 41 660 54
rect 662 45 670 54
rect 662 43 665 45
rect 667 43 670 45
rect 662 41 670 43
rect 620 39 627 41
rect 665 38 670 41
rect 672 38 677 63
rect 679 62 688 63
rect 690 62 695 64
rect 679 57 695 62
rect 679 55 688 57
rect 690 55 695 57
rect 679 38 695 55
rect 697 56 705 66
rect 697 54 700 56
rect 702 54 705 56
rect 697 49 705 54
rect 697 47 700 49
rect 702 47 705 49
rect 697 38 705 47
rect 707 64 715 66
rect 707 62 710 64
rect 712 62 715 64
rect 707 57 715 62
rect 707 55 710 57
rect 712 55 715 57
rect 707 38 715 55
rect 717 51 722 66
rect 732 51 737 66
rect 717 49 724 51
rect 717 47 720 49
rect 722 47 724 49
rect 717 42 724 47
rect 717 40 720 42
rect 722 40 724 42
rect 717 38 724 40
rect 730 49 737 51
rect 730 47 732 49
rect 734 47 737 49
rect 730 42 737 47
rect 730 40 732 42
rect 734 40 737 42
rect 730 38 737 40
rect 739 64 747 66
rect 739 62 742 64
rect 744 62 747 64
rect 739 57 747 62
rect 739 55 742 57
rect 744 55 747 57
rect 739 38 747 55
rect 749 56 757 66
rect 749 54 752 56
rect 754 54 757 56
rect 749 49 757 54
rect 749 47 752 49
rect 754 47 757 49
rect 749 38 757 47
rect 759 64 773 66
rect 759 62 764 64
rect 766 63 773 64
rect 796 64 805 66
rect 766 62 775 63
rect 759 57 775 62
rect 759 55 764 57
rect 766 55 775 57
rect 759 38 775 55
rect 777 38 782 63
rect 784 54 789 63
rect 796 62 799 64
rect 801 62 805 64
rect 796 54 805 62
rect 784 45 792 54
rect 784 43 787 45
rect 789 43 792 45
rect 784 41 792 43
rect 794 41 805 54
rect 807 54 812 66
rect 821 59 826 66
rect 819 57 826 59
rect 819 55 821 57
rect 823 55 826 57
rect 807 52 814 54
rect 819 53 826 55
rect 807 50 810 52
rect 812 50 814 52
rect 807 45 814 50
rect 821 45 826 53
rect 828 45 833 66
rect 835 64 844 66
rect 835 62 840 64
rect 842 62 844 64
rect 835 56 844 62
rect 867 57 874 59
rect 835 45 846 56
rect 807 43 810 45
rect 812 43 814 45
rect 807 41 814 43
rect 784 38 789 41
rect 838 38 846 45
rect 848 54 855 56
rect 848 52 851 54
rect 853 52 855 54
rect 848 47 855 52
rect 848 45 851 47
rect 853 45 855 47
rect 867 55 869 57
rect 871 55 874 57
rect 867 46 874 55
rect 876 57 884 59
rect 876 55 879 57
rect 881 55 884 57
rect 876 50 884 55
rect 876 48 879 50
rect 881 48 884 50
rect 876 46 884 48
rect 886 57 892 59
rect 886 55 894 57
rect 886 53 889 55
rect 891 53 894 55
rect 886 46 894 53
rect 848 43 855 45
rect 848 38 853 43
rect 888 39 894 46
rect 896 52 901 57
rect 919 54 924 66
rect 917 52 924 54
rect 896 50 903 52
rect 896 48 899 50
rect 901 48 903 50
rect 896 43 903 48
rect 896 41 899 43
rect 901 41 903 43
rect 917 50 919 52
rect 921 50 924 52
rect 917 45 924 50
rect 917 43 919 45
rect 921 43 924 45
rect 917 41 924 43
rect 926 64 935 66
rect 926 62 930 64
rect 932 62 935 64
rect 958 64 972 66
rect 958 63 965 64
rect 926 54 935 62
rect 942 54 947 63
rect 926 41 937 54
rect 939 45 947 54
rect 939 43 942 45
rect 944 43 947 45
rect 939 41 947 43
rect 896 39 903 41
rect 942 38 947 41
rect 949 38 954 63
rect 956 62 965 63
rect 967 62 972 64
rect 956 57 972 62
rect 956 55 965 57
rect 967 55 972 57
rect 956 38 972 55
rect 974 56 982 66
rect 974 54 977 56
rect 979 54 982 56
rect 974 49 982 54
rect 974 47 977 49
rect 979 47 982 49
rect 974 38 982 47
rect 984 64 992 66
rect 984 62 987 64
rect 989 62 992 64
rect 984 57 992 62
rect 984 55 987 57
rect 989 55 992 57
rect 984 38 992 55
rect 994 51 999 66
rect 1009 51 1014 66
rect 994 49 1001 51
rect 994 47 997 49
rect 999 47 1001 49
rect 994 42 1001 47
rect 994 40 997 42
rect 999 40 1001 42
rect 994 38 1001 40
rect 1007 49 1014 51
rect 1007 47 1009 49
rect 1011 47 1014 49
rect 1007 42 1014 47
rect 1007 40 1009 42
rect 1011 40 1014 42
rect 1007 38 1014 40
rect 1016 64 1024 66
rect 1016 62 1019 64
rect 1021 62 1024 64
rect 1016 57 1024 62
rect 1016 55 1019 57
rect 1021 55 1024 57
rect 1016 38 1024 55
rect 1026 56 1034 66
rect 1026 54 1029 56
rect 1031 54 1034 56
rect 1026 49 1034 54
rect 1026 47 1029 49
rect 1031 47 1034 49
rect 1026 38 1034 47
rect 1036 64 1050 66
rect 1036 62 1041 64
rect 1043 63 1050 64
rect 1073 64 1082 66
rect 1043 62 1052 63
rect 1036 57 1052 62
rect 1036 55 1041 57
rect 1043 55 1052 57
rect 1036 38 1052 55
rect 1054 38 1059 63
rect 1061 54 1066 63
rect 1073 62 1076 64
rect 1078 62 1082 64
rect 1073 54 1082 62
rect 1061 45 1069 54
rect 1061 43 1064 45
rect 1066 43 1069 45
rect 1061 41 1069 43
rect 1071 41 1082 54
rect 1084 54 1089 66
rect 1098 59 1103 66
rect 1096 57 1103 59
rect 1096 55 1098 57
rect 1100 55 1103 57
rect 1084 52 1091 54
rect 1096 53 1103 55
rect 1084 50 1087 52
rect 1089 50 1091 52
rect 1084 45 1091 50
rect 1098 45 1103 53
rect 1105 45 1110 66
rect 1112 64 1121 66
rect 1112 62 1117 64
rect 1119 62 1121 64
rect 1112 56 1121 62
rect 1112 45 1123 56
rect 1084 43 1087 45
rect 1089 43 1091 45
rect 1084 41 1091 43
rect 1061 38 1066 41
rect 1115 38 1123 45
rect 1125 54 1132 56
rect 1125 52 1128 54
rect 1130 52 1132 54
rect 1125 47 1132 52
rect 1125 45 1128 47
rect 1130 45 1132 47
rect 1125 43 1132 45
rect 1125 38 1130 43
rect -154 -51 -149 -45
rect -156 -53 -149 -51
rect -156 -55 -154 -53
rect -152 -55 -149 -53
rect -156 -57 -149 -55
rect -147 -56 -139 -45
rect -137 -47 -129 -45
rect -137 -49 -134 -47
rect -132 -49 -129 -47
rect -137 -56 -129 -49
rect -127 -46 -119 -45
rect -127 -56 -117 -46
rect -147 -57 -141 -56
rect -145 -62 -141 -57
rect -125 -57 -117 -56
rect -115 -51 -110 -46
rect -102 -51 -97 -45
rect -115 -53 -108 -51
rect -115 -55 -112 -53
rect -110 -55 -108 -53
rect -115 -57 -108 -55
rect -104 -53 -97 -51
rect -104 -55 -102 -53
rect -100 -55 -97 -53
rect -104 -57 -97 -55
rect -95 -56 -87 -45
rect -85 -47 -77 -45
rect -85 -49 -82 -47
rect -80 -49 -77 -47
rect -85 -56 -77 -49
rect -75 -46 -67 -45
rect -75 -56 -65 -46
rect -95 -57 -89 -56
rect -145 -64 -139 -62
rect -145 -66 -143 -64
rect -141 -66 -139 -64
rect -145 -68 -139 -66
rect -125 -64 -119 -57
rect -93 -62 -89 -57
rect -73 -57 -65 -56
rect -63 -51 -58 -46
rect -50 -51 -45 -45
rect -63 -53 -56 -51
rect -63 -55 -60 -53
rect -58 -55 -56 -53
rect -63 -57 -56 -55
rect -52 -53 -45 -51
rect -52 -55 -50 -53
rect -48 -55 -45 -53
rect -52 -57 -45 -55
rect -43 -56 -35 -45
rect -33 -47 -25 -45
rect -33 -49 -30 -47
rect -28 -49 -25 -47
rect -33 -56 -25 -49
rect -23 -46 -15 -45
rect -23 -56 -13 -46
rect -43 -57 -37 -56
rect -125 -66 -123 -64
rect -121 -66 -119 -64
rect -125 -68 -119 -66
rect -93 -64 -87 -62
rect -93 -66 -91 -64
rect -89 -66 -87 -64
rect -93 -68 -87 -66
rect -73 -64 -67 -57
rect -41 -62 -37 -57
rect -21 -57 -13 -56
rect -11 -51 -6 -46
rect 2 -51 7 -45
rect -11 -53 -4 -51
rect -11 -55 -8 -53
rect -6 -55 -4 -53
rect -11 -57 -4 -55
rect 0 -53 7 -51
rect 0 -55 2 -53
rect 4 -55 7 -53
rect 0 -57 7 -55
rect 9 -56 17 -45
rect 19 -47 27 -45
rect 19 -49 22 -47
rect 24 -49 27 -47
rect 19 -56 27 -49
rect 29 -46 37 -45
rect 29 -56 39 -46
rect 9 -57 15 -56
rect -73 -66 -71 -64
rect -69 -66 -67 -64
rect -73 -68 -67 -66
rect -41 -64 -35 -62
rect -41 -66 -39 -64
rect -37 -66 -35 -64
rect -41 -68 -35 -66
rect -21 -64 -15 -57
rect 11 -62 15 -57
rect 31 -57 39 -56
rect 41 -51 46 -46
rect 54 -51 59 -45
rect 41 -53 48 -51
rect 41 -55 44 -53
rect 46 -55 48 -53
rect 41 -57 48 -55
rect 52 -53 59 -51
rect 52 -55 54 -53
rect 56 -55 59 -53
rect 52 -57 59 -55
rect 61 -56 69 -45
rect 71 -47 79 -45
rect 71 -49 74 -47
rect 76 -49 79 -47
rect 71 -56 79 -49
rect 81 -46 89 -45
rect 81 -56 91 -46
rect 61 -57 67 -56
rect -21 -66 -19 -64
rect -17 -66 -15 -64
rect -21 -68 -15 -66
rect 11 -64 17 -62
rect 11 -66 13 -64
rect 15 -66 17 -64
rect 11 -68 17 -66
rect 31 -64 37 -57
rect 63 -62 67 -57
rect 83 -57 91 -56
rect 93 -51 98 -46
rect 107 -51 112 -45
rect 93 -53 100 -51
rect 93 -55 96 -53
rect 98 -55 100 -53
rect 93 -57 100 -55
rect 105 -53 112 -51
rect 105 -55 107 -53
rect 109 -55 112 -53
rect 105 -57 112 -55
rect 114 -56 122 -45
rect 124 -47 132 -45
rect 124 -49 127 -47
rect 129 -49 132 -47
rect 124 -56 132 -49
rect 134 -46 142 -45
rect 134 -56 144 -46
rect 114 -57 120 -56
rect 31 -66 33 -64
rect 35 -66 37 -64
rect 31 -68 37 -66
rect 63 -64 69 -62
rect 63 -66 65 -64
rect 67 -66 69 -64
rect 63 -68 69 -66
rect 83 -64 89 -57
rect 116 -62 120 -57
rect 136 -57 144 -56
rect 146 -51 151 -46
rect 162 -49 169 -37
rect 171 -39 178 -37
rect 171 -41 174 -39
rect 176 -41 178 -39
rect 171 -43 178 -41
rect 171 -49 176 -43
rect 182 -49 189 -37
rect 191 -39 198 -37
rect 191 -41 194 -39
rect 196 -41 198 -39
rect 191 -43 198 -41
rect 191 -49 196 -43
rect 202 -49 209 -37
rect 211 -39 218 -37
rect 211 -41 214 -39
rect 216 -41 218 -39
rect 211 -43 218 -41
rect 211 -49 216 -43
rect 224 -49 231 -37
rect 233 -39 240 -37
rect 233 -41 236 -39
rect 238 -41 240 -39
rect 233 -43 240 -41
rect 233 -49 238 -43
rect 246 -49 253 -37
rect 255 -39 262 -37
rect 255 -41 258 -39
rect 260 -41 262 -39
rect 255 -43 262 -41
rect 255 -49 260 -43
rect 268 -49 275 -37
rect 277 -39 284 -37
rect 277 -41 280 -39
rect 282 -41 284 -39
rect 277 -43 284 -41
rect 277 -49 282 -43
rect 146 -53 153 -51
rect 146 -55 149 -53
rect 151 -55 153 -53
rect 146 -57 153 -55
rect 83 -66 85 -64
rect 87 -66 89 -64
rect 83 -68 89 -66
rect 116 -64 122 -62
rect 116 -66 118 -64
rect 120 -66 122 -64
rect 116 -68 122 -66
rect 136 -64 142 -57
rect 162 -60 167 -49
rect 182 -60 187 -49
rect 202 -60 207 -49
rect 224 -60 229 -49
rect 246 -60 251 -49
rect 268 -60 273 -49
rect 295 -51 300 -45
rect 293 -53 300 -51
rect 293 -55 295 -53
rect 297 -55 300 -53
rect 293 -57 300 -55
rect 302 -56 310 -45
rect 312 -47 320 -45
rect 312 -49 315 -47
rect 317 -49 320 -47
rect 312 -56 320 -49
rect 322 -46 330 -45
rect 322 -56 332 -46
rect 302 -57 308 -56
rect 136 -66 138 -64
rect 140 -66 142 -64
rect 136 -68 142 -66
rect 162 -64 168 -60
rect 162 -66 164 -64
rect 166 -66 168 -64
rect 162 -68 168 -66
rect 182 -64 188 -60
rect 182 -66 184 -64
rect 186 -66 188 -64
rect 182 -68 188 -66
rect 202 -64 208 -60
rect 202 -66 204 -64
rect 206 -66 208 -64
rect 202 -68 208 -66
rect 224 -64 230 -60
rect 224 -66 226 -64
rect 228 -66 230 -64
rect 224 -68 230 -66
rect 246 -64 252 -60
rect 246 -66 248 -64
rect 250 -66 252 -64
rect 246 -68 252 -66
rect 268 -64 274 -60
rect 268 -66 270 -64
rect 272 -66 274 -64
rect 268 -68 274 -66
rect 304 -62 308 -57
rect 324 -57 332 -56
rect 334 -51 339 -46
rect 348 -51 353 -45
rect 334 -53 341 -51
rect 334 -55 337 -53
rect 339 -55 341 -53
rect 334 -57 341 -55
rect 346 -53 353 -51
rect 346 -55 348 -53
rect 350 -55 353 -53
rect 346 -57 353 -55
rect 355 -56 363 -45
rect 365 -47 373 -45
rect 365 -49 368 -47
rect 370 -49 373 -47
rect 365 -56 373 -49
rect 375 -46 383 -45
rect 375 -56 385 -46
rect 355 -57 361 -56
rect 304 -64 310 -62
rect 304 -66 306 -64
rect 308 -66 310 -64
rect 304 -68 310 -66
rect 324 -64 330 -57
rect 357 -62 361 -57
rect 377 -57 385 -56
rect 387 -51 392 -46
rect 400 -51 405 -45
rect 387 -53 394 -51
rect 387 -55 390 -53
rect 392 -55 394 -53
rect 387 -57 394 -55
rect 398 -53 405 -51
rect 398 -55 400 -53
rect 402 -55 405 -53
rect 398 -57 405 -55
rect 407 -56 415 -45
rect 417 -47 425 -45
rect 417 -49 420 -47
rect 422 -49 425 -47
rect 417 -56 425 -49
rect 427 -46 435 -45
rect 427 -56 437 -46
rect 407 -57 413 -56
rect 324 -66 326 -64
rect 328 -66 330 -64
rect 324 -68 330 -66
rect 357 -64 363 -62
rect 357 -66 359 -64
rect 361 -66 363 -64
rect 357 -68 363 -66
rect 377 -64 383 -57
rect 409 -62 413 -57
rect 429 -57 437 -56
rect 439 -51 444 -46
rect 452 -51 457 -45
rect 439 -53 446 -51
rect 439 -55 442 -53
rect 444 -55 446 -53
rect 439 -57 446 -55
rect 450 -53 457 -51
rect 450 -55 452 -53
rect 454 -55 457 -53
rect 450 -57 457 -55
rect 459 -56 467 -45
rect 469 -47 477 -45
rect 469 -49 472 -47
rect 474 -49 477 -47
rect 469 -56 477 -49
rect 479 -46 487 -45
rect 479 -56 489 -46
rect 459 -57 465 -56
rect 377 -66 379 -64
rect 381 -66 383 -64
rect 377 -68 383 -66
rect 409 -64 415 -62
rect 409 -66 411 -64
rect 413 -66 415 -64
rect 409 -68 415 -66
rect 429 -64 435 -57
rect 461 -62 465 -57
rect 481 -57 489 -56
rect 491 -51 496 -46
rect 504 -51 509 -45
rect 491 -53 498 -51
rect 491 -55 494 -53
rect 496 -55 498 -53
rect 491 -57 498 -55
rect 502 -53 509 -51
rect 502 -55 504 -53
rect 506 -55 509 -53
rect 502 -57 509 -55
rect 511 -56 519 -45
rect 521 -47 529 -45
rect 521 -49 524 -47
rect 526 -49 529 -47
rect 521 -56 529 -49
rect 531 -46 539 -45
rect 531 -56 541 -46
rect 511 -57 517 -56
rect 429 -66 431 -64
rect 433 -66 435 -64
rect 429 -68 435 -66
rect 461 -64 467 -62
rect 461 -66 463 -64
rect 465 -66 467 -64
rect 461 -68 467 -66
rect 481 -64 487 -57
rect 513 -62 517 -57
rect 533 -57 541 -56
rect 543 -51 548 -46
rect 557 -49 564 -37
rect 566 -39 573 -37
rect 566 -41 569 -39
rect 571 -41 573 -39
rect 566 -43 573 -41
rect 566 -49 571 -43
rect 578 -49 585 -37
rect 587 -39 594 -37
rect 587 -41 590 -39
rect 592 -41 594 -39
rect 587 -43 594 -41
rect 587 -49 592 -43
rect 543 -53 550 -51
rect 543 -55 546 -53
rect 548 -55 550 -53
rect 543 -57 550 -55
rect 481 -66 483 -64
rect 485 -66 487 -64
rect 481 -68 487 -66
rect 513 -64 519 -62
rect 513 -66 515 -64
rect 517 -66 519 -64
rect 513 -68 519 -66
rect 533 -64 539 -57
rect 557 -60 562 -49
rect 578 -60 583 -49
rect 603 -51 608 -45
rect 601 -53 608 -51
rect 601 -55 603 -53
rect 605 -55 608 -53
rect 601 -57 608 -55
rect 610 -56 618 -45
rect 620 -47 628 -45
rect 620 -49 623 -47
rect 625 -49 628 -47
rect 620 -56 628 -49
rect 630 -46 638 -45
rect 630 -56 640 -46
rect 610 -57 616 -56
rect 533 -66 535 -64
rect 537 -66 539 -64
rect 533 -68 539 -66
rect 557 -64 563 -60
rect 557 -66 559 -64
rect 561 -66 563 -64
rect 557 -68 563 -66
rect 578 -64 584 -60
rect 578 -66 580 -64
rect 582 -66 584 -64
rect 578 -68 584 -66
rect 612 -62 616 -57
rect 632 -57 640 -56
rect 642 -51 647 -46
rect 656 -51 661 -45
rect 642 -53 649 -51
rect 642 -55 645 -53
rect 647 -55 649 -53
rect 642 -57 649 -55
rect 654 -53 661 -51
rect 654 -55 656 -53
rect 658 -55 661 -53
rect 654 -57 661 -55
rect 663 -56 671 -45
rect 673 -47 681 -45
rect 673 -49 676 -47
rect 678 -49 681 -47
rect 673 -56 681 -49
rect 683 -46 691 -45
rect 683 -56 693 -46
rect 663 -57 669 -56
rect 612 -64 618 -62
rect 612 -66 614 -64
rect 616 -66 618 -64
rect 612 -68 618 -66
rect 632 -64 638 -57
rect 665 -62 669 -57
rect 685 -57 693 -56
rect 695 -51 700 -46
rect 708 -51 713 -45
rect 695 -53 702 -51
rect 695 -55 698 -53
rect 700 -55 702 -53
rect 695 -57 702 -55
rect 706 -53 713 -51
rect 706 -55 708 -53
rect 710 -55 713 -53
rect 706 -57 713 -55
rect 715 -56 723 -45
rect 725 -47 733 -45
rect 725 -49 728 -47
rect 730 -49 733 -47
rect 725 -56 733 -49
rect 735 -46 743 -45
rect 735 -56 745 -46
rect 715 -57 721 -56
rect 632 -66 634 -64
rect 636 -66 638 -64
rect 632 -68 638 -66
rect 665 -64 671 -62
rect 665 -66 667 -64
rect 669 -66 671 -64
rect 665 -68 671 -66
rect 685 -64 691 -57
rect 717 -62 721 -57
rect 737 -57 745 -56
rect 747 -51 752 -46
rect 760 -51 765 -45
rect 747 -53 754 -51
rect 747 -55 750 -53
rect 752 -55 754 -53
rect 747 -57 754 -55
rect 758 -53 765 -51
rect 758 -55 760 -53
rect 762 -55 765 -53
rect 758 -57 765 -55
rect 767 -56 775 -45
rect 777 -47 785 -45
rect 777 -49 780 -47
rect 782 -49 785 -47
rect 777 -56 785 -49
rect 787 -46 795 -45
rect 787 -56 797 -46
rect 767 -57 773 -56
rect 685 -66 687 -64
rect 689 -66 691 -64
rect 685 -68 691 -66
rect 717 -64 723 -62
rect 717 -66 719 -64
rect 721 -66 723 -64
rect 717 -68 723 -66
rect 737 -64 743 -57
rect 769 -62 773 -57
rect 789 -57 797 -56
rect 799 -51 804 -46
rect 812 -51 817 -45
rect 799 -53 806 -51
rect 799 -55 802 -53
rect 804 -55 806 -53
rect 799 -57 806 -55
rect 810 -53 817 -51
rect 810 -55 812 -53
rect 814 -55 817 -53
rect 810 -57 817 -55
rect 819 -56 827 -45
rect 829 -47 837 -45
rect 829 -49 832 -47
rect 834 -49 837 -47
rect 829 -56 837 -49
rect 839 -46 847 -45
rect 839 -56 849 -46
rect 819 -57 825 -56
rect 737 -66 739 -64
rect 741 -66 743 -64
rect 737 -68 743 -66
rect 769 -64 775 -62
rect 769 -66 771 -64
rect 773 -66 775 -64
rect 769 -68 775 -66
rect 789 -64 795 -57
rect 821 -62 825 -57
rect 841 -57 849 -56
rect 851 -51 856 -46
rect 864 -51 869 -45
rect 851 -53 858 -51
rect 851 -55 854 -53
rect 856 -55 858 -53
rect 851 -57 858 -55
rect 862 -53 869 -51
rect 862 -55 864 -53
rect 866 -55 869 -53
rect 862 -57 869 -55
rect 871 -56 879 -45
rect 881 -47 889 -45
rect 881 -49 884 -47
rect 886 -49 889 -47
rect 881 -56 889 -49
rect 891 -46 899 -45
rect 891 -56 901 -46
rect 871 -57 877 -56
rect 789 -66 791 -64
rect 793 -66 795 -64
rect 789 -68 795 -66
rect 821 -64 827 -62
rect 821 -66 823 -64
rect 825 -66 827 -64
rect 821 -68 827 -66
rect 841 -64 847 -57
rect 873 -62 877 -57
rect 893 -57 901 -56
rect 903 -51 908 -46
rect 917 -51 922 -45
rect 903 -53 910 -51
rect 903 -55 906 -53
rect 908 -55 910 -53
rect 903 -57 910 -55
rect 915 -53 922 -51
rect 915 -55 917 -53
rect 919 -55 922 -53
rect 915 -57 922 -55
rect 924 -56 932 -45
rect 934 -47 942 -45
rect 934 -49 937 -47
rect 939 -49 942 -47
rect 934 -56 942 -49
rect 944 -46 952 -45
rect 944 -56 954 -46
rect 924 -57 930 -56
rect 841 -66 843 -64
rect 845 -66 847 -64
rect 841 -68 847 -66
rect 873 -64 879 -62
rect 873 -66 875 -64
rect 877 -66 879 -64
rect 873 -68 879 -66
rect 893 -64 899 -57
rect 926 -62 930 -57
rect 946 -57 954 -56
rect 956 -51 961 -46
rect 971 -51 976 -45
rect 956 -53 963 -51
rect 956 -55 959 -53
rect 961 -55 963 -53
rect 956 -57 963 -55
rect 969 -53 976 -51
rect 969 -55 971 -53
rect 973 -55 976 -53
rect 969 -57 976 -55
rect 978 -56 986 -45
rect 988 -47 996 -45
rect 988 -49 991 -47
rect 993 -49 996 -47
rect 988 -56 996 -49
rect 998 -46 1006 -45
rect 998 -56 1008 -46
rect 978 -57 984 -56
rect 893 -66 895 -64
rect 897 -66 899 -64
rect 893 -68 899 -66
rect 926 -64 932 -62
rect 926 -66 928 -64
rect 930 -66 932 -64
rect 926 -68 932 -66
rect 946 -64 952 -57
rect 980 -62 984 -57
rect 1000 -57 1008 -56
rect 1010 -51 1015 -46
rect 1026 -51 1031 -45
rect 1010 -53 1017 -51
rect 1010 -55 1013 -53
rect 1015 -55 1017 -53
rect 1010 -57 1017 -55
rect 1024 -53 1031 -51
rect 1024 -55 1026 -53
rect 1028 -55 1031 -53
rect 1024 -57 1031 -55
rect 1033 -56 1041 -45
rect 1043 -47 1051 -45
rect 1043 -49 1046 -47
rect 1048 -49 1051 -47
rect 1043 -56 1051 -49
rect 1053 -46 1061 -45
rect 1053 -56 1063 -46
rect 1033 -57 1039 -56
rect 946 -66 948 -64
rect 950 -66 952 -64
rect 946 -68 952 -66
rect 980 -64 986 -62
rect 980 -66 982 -64
rect 984 -66 986 -64
rect 980 -68 986 -66
rect 1000 -64 1006 -57
rect 1035 -62 1039 -57
rect 1055 -57 1063 -56
rect 1065 -51 1070 -46
rect 1079 -51 1084 -45
rect 1065 -53 1072 -51
rect 1065 -55 1068 -53
rect 1070 -55 1072 -53
rect 1065 -57 1072 -55
rect 1077 -53 1084 -51
rect 1077 -55 1079 -53
rect 1081 -55 1084 -53
rect 1077 -57 1084 -55
rect 1086 -56 1094 -45
rect 1096 -47 1104 -45
rect 1096 -49 1099 -47
rect 1101 -49 1104 -47
rect 1096 -56 1104 -49
rect 1106 -46 1114 -45
rect 1106 -56 1116 -46
rect 1086 -57 1092 -56
rect 1000 -66 1002 -64
rect 1004 -66 1006 -64
rect 1000 -68 1006 -66
rect 1035 -64 1041 -62
rect 1035 -66 1037 -64
rect 1039 -66 1041 -64
rect 1035 -68 1041 -66
rect 1055 -64 1061 -57
rect 1088 -62 1092 -57
rect 1108 -57 1116 -56
rect 1118 -51 1123 -46
rect 1118 -53 1125 -51
rect 1118 -55 1121 -53
rect 1123 -55 1125 -53
rect 1118 -57 1125 -55
rect 1055 -66 1057 -64
rect 1059 -66 1061 -64
rect 1055 -68 1061 -66
rect 1088 -64 1094 -62
rect 1088 -66 1090 -64
rect 1092 -66 1094 -64
rect 1088 -68 1094 -66
rect 1108 -64 1114 -57
rect 1108 -66 1110 -64
rect 1112 -66 1114 -64
rect 1108 -68 1114 -66
<< alu1 >>
rect -290 358 1136 360
rect -290 356 98 358
rect 100 356 1136 358
rect -290 355 1136 356
rect -290 353 -247 355
rect -245 353 -5 355
rect -3 353 38 355
rect 40 353 78 355
rect 80 353 297 355
rect 299 353 345 355
rect 347 353 574 355
rect 576 353 622 355
rect 624 353 850 355
rect 852 353 898 355
rect 900 353 1127 355
rect 1129 353 1136 355
rect -290 352 1136 353
rect -283 344 -271 347
rect -283 342 -276 344
rect -274 342 -271 344
rect -290 341 -271 342
rect -290 338 -278 341
rect -283 329 -278 338
rect -4 346 0 347
rect -13 342 0 346
rect -215 340 -210 342
rect -283 327 -281 329
rect -279 327 -278 329
rect -283 325 -278 327
rect -267 322 -262 323
rect -267 320 -265 322
rect -263 320 -262 322
rect -267 316 -262 320
rect -239 338 -223 339
rect -239 336 -237 338
rect -235 336 -223 338
rect -239 334 -223 336
rect -227 322 -223 334
rect -227 320 -226 322
rect -224 320 -223 322
rect -267 315 -265 316
rect -275 314 -265 315
rect -263 314 -262 316
rect -275 313 -262 314
rect -275 311 -274 313
rect -272 312 -262 313
rect -272 311 -265 312
rect -275 310 -265 311
rect -263 310 -262 312
rect -275 309 -262 310
rect -227 306 -223 320
rect -247 305 -223 306
rect -247 303 -245 305
rect -243 303 -223 305
rect -247 302 -223 303
rect -215 338 -213 340
rect -211 338 -210 340
rect -215 333 -210 338
rect -215 331 -213 333
rect -211 331 -210 333
rect -215 329 -210 331
rect -215 313 -211 329
rect -184 326 -146 330
rect -184 323 -179 326
rect -187 322 -179 323
rect -187 321 -182 322
rect -187 319 -186 321
rect -184 320 -182 321
rect -180 320 -179 322
rect -184 319 -179 320
rect -187 317 -179 319
rect -169 321 -154 322
rect -169 319 -167 321
rect -165 319 -160 321
rect -158 319 -157 321
rect -155 319 -154 321
rect -169 318 -154 319
rect -215 311 -214 313
rect -212 311 -211 313
rect -215 307 -211 311
rect -215 305 -210 307
rect -167 309 -163 318
rect -136 337 -130 339
rect -136 335 -135 337
rect -133 335 -130 337
rect -136 330 -130 335
rect -136 328 -135 330
rect -133 328 -130 330
rect -136 326 -130 328
rect -134 321 -130 326
rect -134 319 -133 321
rect -131 319 -130 321
rect -134 306 -130 319
rect -215 303 -213 305
rect -211 303 -210 305
rect -215 301 -210 303
rect -136 305 -130 306
rect -136 303 -135 305
rect -133 303 -130 305
rect -136 302 -130 303
rect -126 337 -120 339
rect -46 340 -41 342
rect -46 338 -45 340
rect -43 338 -41 340
rect -126 335 -123 337
rect -121 335 -120 337
rect -126 334 -120 335
rect -126 332 -123 334
rect -121 332 -120 334
rect -126 330 -120 332
rect -126 328 -123 330
rect -121 328 -120 330
rect -126 326 -120 328
rect -126 306 -122 326
rect -110 329 -72 330
rect -110 327 -104 329
rect -102 327 -72 329
rect -110 326 -72 327
rect -77 323 -72 326
rect -102 321 -87 322
rect -102 319 -98 321
rect -96 319 -91 321
rect -89 319 -87 321
rect -102 318 -87 319
rect -77 321 -69 323
rect -77 319 -72 321
rect -70 319 -69 321
rect -93 313 -89 318
rect -77 317 -69 319
rect -46 333 -41 338
rect -46 331 -45 333
rect -43 331 -41 333
rect -46 329 -41 331
rect -93 311 -92 313
rect -90 311 -89 313
rect -93 309 -89 311
rect -126 305 -120 306
rect -126 303 -123 305
rect -121 303 -120 305
rect -126 302 -120 303
rect -45 309 -41 329
rect -36 334 -32 339
rect -36 332 -35 334
rect -33 332 -32 334
rect -36 330 -32 332
rect -36 328 -15 330
rect -36 326 -31 328
rect -29 326 -15 328
rect -36 321 -15 322
rect -36 319 -35 321
rect -33 319 -21 321
rect -19 319 -15 321
rect -36 318 -15 319
rect -2 340 0 342
rect -4 335 0 340
rect -2 333 0 335
rect -36 309 -32 318
rect -4 317 0 333
rect 7 332 11 339
rect 38 338 43 340
rect 7 330 8 332
rect 10 330 11 332
rect 7 329 20 330
rect 7 327 12 329
rect 14 327 20 329
rect 7 326 20 327
rect -4 315 -3 317
rect -1 315 0 317
rect -4 314 0 315
rect -5 312 0 314
rect -5 310 -4 312
rect -2 310 0 312
rect -45 307 -44 309
rect -42 307 -41 309
rect -5 308 0 310
rect 14 321 28 322
rect 14 319 22 321
rect 24 319 28 321
rect 14 318 28 319
rect 38 336 39 338
rect 41 336 43 338
rect 38 331 43 336
rect 38 329 39 331
rect 41 329 43 331
rect 38 327 43 329
rect 14 312 19 318
rect 14 310 16 312
rect 18 310 19 312
rect 14 309 19 310
rect 39 326 43 327
rect 47 338 51 339
rect 47 336 48 338
rect 50 336 51 338
rect 47 330 51 336
rect 298 346 302 347
rect 289 342 302 346
rect 87 340 92 342
rect 78 338 83 340
rect 47 329 60 330
rect 47 327 52 329
rect 54 327 60 329
rect 47 326 60 327
rect 39 324 40 326
rect 42 324 43 326
rect -46 305 -41 307
rect 39 307 43 324
rect 54 321 68 322
rect 54 319 62 321
rect 64 319 68 321
rect 54 318 68 319
rect 78 336 79 338
rect 81 336 83 338
rect 78 331 83 336
rect 78 329 79 331
rect 81 329 83 331
rect 78 327 83 329
rect 54 315 59 318
rect 54 313 56 315
rect 58 313 59 315
rect 54 309 59 313
rect 79 321 83 327
rect 79 319 80 321
rect 82 319 83 321
rect -46 303 -45 305
rect -43 303 -41 305
rect -46 301 -41 303
rect 31 305 39 307
rect 41 305 43 307
rect 79 307 83 319
rect 31 301 43 305
rect 71 305 79 307
rect 81 305 83 307
rect 71 301 83 305
rect 87 338 89 340
rect 91 338 92 340
rect 87 333 92 338
rect 87 331 89 333
rect 91 331 92 333
rect 87 329 92 331
rect 87 313 91 329
rect 118 329 156 330
rect 118 327 120 329
rect 122 327 156 329
rect 118 326 156 327
rect 118 323 123 326
rect 115 321 123 323
rect 115 319 116 321
rect 118 319 123 321
rect 115 317 123 319
rect 133 321 148 322
rect 133 319 135 321
rect 137 319 138 321
rect 140 319 142 321
rect 144 319 148 321
rect 133 318 148 319
rect 87 311 88 313
rect 90 311 91 313
rect 87 307 91 311
rect 87 305 92 307
rect 135 309 139 318
rect 166 337 172 339
rect 166 335 167 337
rect 169 335 172 337
rect 166 330 172 335
rect 166 328 167 330
rect 169 328 172 330
rect 166 326 172 328
rect 168 321 172 326
rect 168 319 169 321
rect 171 319 172 321
rect 168 306 172 319
rect 87 303 89 305
rect 91 303 92 305
rect 87 301 92 303
rect 166 305 172 306
rect 166 303 167 305
rect 169 303 172 305
rect 166 302 172 303
rect 176 337 182 339
rect 256 340 261 342
rect 256 338 257 340
rect 259 338 261 340
rect 176 335 179 337
rect 181 335 182 337
rect 176 334 182 335
rect 176 332 179 334
rect 181 332 182 334
rect 176 330 182 332
rect 176 328 179 330
rect 181 328 182 330
rect 176 326 182 328
rect 176 306 180 326
rect 192 329 230 330
rect 192 327 209 329
rect 211 327 230 329
rect 192 326 230 327
rect 225 323 230 326
rect 200 321 215 322
rect 200 319 204 321
rect 206 319 211 321
rect 213 319 215 321
rect 200 318 215 319
rect 225 321 233 323
rect 225 319 230 321
rect 232 319 233 321
rect 209 313 213 318
rect 225 317 233 319
rect 256 333 261 338
rect 256 331 257 333
rect 259 331 261 333
rect 256 329 261 331
rect 209 311 210 313
rect 212 311 213 313
rect 209 309 213 311
rect 176 305 182 306
rect 176 303 179 305
rect 181 303 182 305
rect 176 302 182 303
rect 257 309 261 329
rect 266 338 270 339
rect 266 336 267 338
rect 269 336 270 338
rect 266 330 270 336
rect 266 328 287 330
rect 266 326 271 328
rect 273 326 287 328
rect 266 321 287 322
rect 266 319 267 321
rect 269 319 281 321
rect 283 319 287 321
rect 266 318 287 319
rect 300 340 302 342
rect 298 335 302 340
rect 300 333 302 335
rect 266 309 270 318
rect 298 317 302 333
rect 314 334 318 339
rect 314 332 315 334
rect 317 332 318 334
rect 575 346 579 347
rect 566 342 579 346
rect 364 340 369 342
rect 345 338 350 340
rect 314 330 318 332
rect 314 329 327 330
rect 314 327 319 329
rect 321 327 327 329
rect 314 326 327 327
rect 298 315 299 317
rect 301 315 302 317
rect 298 314 302 315
rect 297 312 302 314
rect 297 310 298 312
rect 300 310 302 312
rect 257 307 258 309
rect 260 307 261 309
rect 297 308 302 310
rect 321 321 335 322
rect 321 319 329 321
rect 331 319 332 321
rect 334 319 335 321
rect 321 318 335 319
rect 345 336 346 338
rect 348 336 350 338
rect 345 331 350 336
rect 345 329 346 331
rect 348 329 350 331
rect 345 327 350 329
rect 321 309 326 318
rect 346 326 350 327
rect 346 324 347 326
rect 349 324 350 326
rect 256 305 261 307
rect 346 307 350 324
rect 256 303 257 305
rect 259 303 261 305
rect 256 301 261 303
rect 338 305 346 307
rect 348 305 350 307
rect 338 301 350 305
rect 364 338 366 340
rect 368 338 369 340
rect 364 333 369 338
rect 364 331 366 333
rect 368 331 369 333
rect 364 329 369 331
rect 364 313 368 329
rect 395 329 433 330
rect 395 327 397 329
rect 399 327 433 329
rect 395 326 433 327
rect 395 323 400 326
rect 392 321 400 323
rect 392 319 393 321
rect 395 319 400 321
rect 392 317 400 319
rect 410 321 425 322
rect 410 319 412 321
rect 414 319 415 321
rect 417 319 419 321
rect 421 319 425 321
rect 410 318 425 319
rect 364 311 365 313
rect 367 311 368 313
rect 364 307 368 311
rect 364 305 369 307
rect 412 309 416 318
rect 443 337 449 339
rect 443 335 444 337
rect 446 335 449 337
rect 443 330 449 335
rect 443 328 444 330
rect 446 328 449 330
rect 443 326 449 328
rect 445 321 449 326
rect 445 319 446 321
rect 448 319 449 321
rect 445 306 449 319
rect 364 303 366 305
rect 368 303 369 305
rect 364 301 369 303
rect 443 305 449 306
rect 443 303 444 305
rect 446 303 449 305
rect 443 302 449 303
rect 453 337 459 339
rect 533 340 538 342
rect 533 338 534 340
rect 536 338 538 340
rect 453 335 456 337
rect 458 335 459 337
rect 453 334 459 335
rect 453 332 456 334
rect 458 332 459 334
rect 453 330 459 332
rect 453 328 456 330
rect 458 328 459 330
rect 453 326 459 328
rect 453 306 457 326
rect 469 329 507 330
rect 469 327 486 329
rect 488 327 507 329
rect 469 326 507 327
rect 502 323 507 326
rect 477 321 492 322
rect 477 319 481 321
rect 483 319 488 321
rect 490 319 492 321
rect 477 318 492 319
rect 502 321 510 323
rect 502 319 507 321
rect 509 319 510 321
rect 486 313 490 318
rect 502 317 510 319
rect 533 333 538 338
rect 533 331 534 333
rect 536 331 538 333
rect 533 329 538 331
rect 486 311 487 313
rect 489 311 490 313
rect 486 309 490 311
rect 453 305 459 306
rect 453 303 456 305
rect 458 303 459 305
rect 453 302 459 303
rect 534 309 538 329
rect 543 338 547 339
rect 543 336 544 338
rect 546 336 547 338
rect 543 330 547 336
rect 543 328 564 330
rect 543 326 548 328
rect 550 326 564 328
rect 543 321 564 322
rect 543 319 544 321
rect 546 319 558 321
rect 560 319 564 321
rect 543 318 564 319
rect 577 340 579 342
rect 575 335 579 340
rect 577 333 579 335
rect 543 309 547 318
rect 575 317 579 333
rect 591 334 595 339
rect 591 332 592 334
rect 594 332 595 334
rect 851 346 855 347
rect 842 342 855 346
rect 640 340 645 342
rect 622 338 627 340
rect 591 330 595 332
rect 591 329 604 330
rect 591 327 596 329
rect 598 327 604 329
rect 591 326 604 327
rect 575 315 576 317
rect 578 315 579 317
rect 575 314 579 315
rect 574 312 579 314
rect 574 310 575 312
rect 577 310 579 312
rect 534 307 535 309
rect 537 307 538 309
rect 574 308 579 310
rect 598 321 612 322
rect 598 319 606 321
rect 608 319 609 321
rect 611 319 612 321
rect 598 318 612 319
rect 622 336 623 338
rect 625 336 627 338
rect 622 331 627 336
rect 622 329 623 331
rect 625 329 627 331
rect 622 327 627 329
rect 598 309 603 318
rect 623 326 627 327
rect 623 324 624 326
rect 626 324 627 326
rect 533 305 538 307
rect 623 307 627 324
rect 533 303 534 305
rect 536 303 538 305
rect 533 301 538 303
rect 615 305 623 307
rect 625 305 627 307
rect 615 301 627 305
rect 640 338 642 340
rect 644 338 645 340
rect 640 333 645 338
rect 640 331 642 333
rect 644 331 645 333
rect 640 329 645 331
rect 640 313 644 329
rect 671 329 709 330
rect 671 327 673 329
rect 675 327 709 329
rect 671 326 709 327
rect 671 323 676 326
rect 668 321 676 323
rect 668 319 669 321
rect 671 319 676 321
rect 668 317 676 319
rect 686 321 701 322
rect 686 319 688 321
rect 690 319 691 321
rect 693 319 695 321
rect 697 319 701 321
rect 686 318 701 319
rect 640 311 641 313
rect 643 311 644 313
rect 640 307 644 311
rect 640 305 645 307
rect 688 309 692 318
rect 719 337 725 339
rect 719 335 720 337
rect 722 335 725 337
rect 719 330 725 335
rect 719 328 720 330
rect 722 328 725 330
rect 719 326 725 328
rect 721 321 725 326
rect 721 319 722 321
rect 724 319 725 321
rect 721 306 725 319
rect 640 303 642 305
rect 644 303 645 305
rect 640 301 645 303
rect 719 305 725 306
rect 719 303 720 305
rect 722 303 725 305
rect 719 302 725 303
rect 729 337 735 339
rect 809 340 814 342
rect 809 338 810 340
rect 812 338 814 340
rect 729 335 732 337
rect 734 335 735 337
rect 729 334 735 335
rect 729 332 732 334
rect 734 332 735 334
rect 729 330 735 332
rect 729 328 732 330
rect 734 328 735 330
rect 729 326 735 328
rect 729 306 733 326
rect 745 329 783 330
rect 745 327 762 329
rect 764 327 783 329
rect 745 326 783 327
rect 778 323 783 326
rect 753 321 768 322
rect 753 319 757 321
rect 759 319 764 321
rect 766 319 768 321
rect 753 318 768 319
rect 778 321 786 323
rect 778 319 783 321
rect 785 319 786 321
rect 762 313 766 318
rect 778 317 786 319
rect 809 333 814 338
rect 809 331 810 333
rect 812 331 814 333
rect 809 329 814 331
rect 762 311 763 313
rect 765 311 766 313
rect 762 309 766 311
rect 729 305 735 306
rect 729 303 732 305
rect 734 303 735 305
rect 729 302 735 303
rect 810 310 814 329
rect 819 338 823 339
rect 819 336 820 338
rect 822 336 823 338
rect 819 330 823 336
rect 819 328 840 330
rect 819 326 824 328
rect 826 326 840 328
rect 810 308 811 310
rect 813 308 814 310
rect 819 321 840 322
rect 819 319 820 321
rect 822 319 834 321
rect 836 319 840 321
rect 819 318 840 319
rect 853 340 855 342
rect 851 335 855 340
rect 853 333 855 335
rect 819 309 823 318
rect 851 317 855 333
rect 867 334 871 339
rect 867 332 868 334
rect 870 332 871 334
rect 1128 346 1132 347
rect 1119 342 1132 346
rect 917 340 922 342
rect 898 338 903 340
rect 867 330 871 332
rect 867 329 880 330
rect 867 327 872 329
rect 874 327 880 329
rect 867 326 880 327
rect 851 315 852 317
rect 854 315 855 317
rect 851 314 855 315
rect 850 312 855 314
rect 850 310 851 312
rect 853 310 855 312
rect 850 308 855 310
rect 874 321 888 322
rect 874 319 882 321
rect 884 319 885 321
rect 887 319 888 321
rect 874 318 888 319
rect 898 336 899 338
rect 901 336 903 338
rect 898 331 903 336
rect 898 329 899 331
rect 901 329 903 331
rect 898 327 903 329
rect 874 309 879 318
rect 899 326 903 327
rect 899 324 900 326
rect 902 324 903 326
rect 810 307 814 308
rect 809 305 814 307
rect 899 307 903 324
rect 809 303 810 305
rect 812 303 814 305
rect 809 301 814 303
rect 891 305 899 307
rect 901 305 903 307
rect 891 301 903 305
rect 917 338 919 340
rect 921 338 922 340
rect 917 333 922 338
rect 917 331 919 333
rect 921 331 922 333
rect 917 329 922 331
rect 917 313 921 329
rect 948 329 986 330
rect 948 327 950 329
rect 952 327 986 329
rect 948 326 986 327
rect 948 323 953 326
rect 945 321 953 323
rect 945 319 946 321
rect 948 319 953 321
rect 945 317 953 319
rect 963 321 978 322
rect 963 319 965 321
rect 967 319 968 321
rect 970 319 972 321
rect 974 319 978 321
rect 963 318 978 319
rect 917 311 918 313
rect 920 311 921 313
rect 917 307 921 311
rect 917 305 922 307
rect 965 309 969 318
rect 996 337 1002 339
rect 996 335 997 337
rect 999 335 1002 337
rect 996 330 1002 335
rect 996 328 997 330
rect 999 328 1002 330
rect 996 326 1002 328
rect 998 321 1002 326
rect 998 319 999 321
rect 1001 319 1002 321
rect 998 306 1002 319
rect 917 303 919 305
rect 921 303 922 305
rect 917 301 922 303
rect 996 305 1002 306
rect 996 303 997 305
rect 999 303 1002 305
rect 996 302 1002 303
rect 1006 337 1012 339
rect 1086 340 1091 342
rect 1086 338 1087 340
rect 1089 338 1091 340
rect 1006 335 1009 337
rect 1011 335 1012 337
rect 1006 334 1012 335
rect 1006 332 1009 334
rect 1011 332 1012 334
rect 1006 330 1012 332
rect 1006 328 1009 330
rect 1011 328 1012 330
rect 1006 326 1012 328
rect 1006 306 1010 326
rect 1022 329 1060 330
rect 1022 327 1039 329
rect 1041 327 1060 329
rect 1022 326 1060 327
rect 1055 323 1060 326
rect 1030 321 1045 322
rect 1030 319 1034 321
rect 1036 319 1041 321
rect 1043 319 1045 321
rect 1030 318 1045 319
rect 1055 321 1063 323
rect 1055 319 1060 321
rect 1062 319 1063 321
rect 1039 313 1043 318
rect 1055 317 1063 319
rect 1086 333 1091 338
rect 1086 331 1087 333
rect 1089 331 1091 333
rect 1086 329 1091 331
rect 1039 311 1040 313
rect 1042 311 1043 313
rect 1039 309 1043 311
rect 1006 305 1012 306
rect 1006 303 1009 305
rect 1011 303 1012 305
rect 1006 302 1012 303
rect 1087 308 1091 329
rect 1096 338 1100 339
rect 1096 336 1097 338
rect 1099 336 1100 338
rect 1096 330 1100 336
rect 1096 328 1117 330
rect 1096 326 1101 328
rect 1103 326 1117 328
rect 1096 321 1117 322
rect 1096 319 1097 321
rect 1099 319 1111 321
rect 1113 319 1117 321
rect 1096 318 1117 319
rect 1130 340 1132 342
rect 1128 335 1132 340
rect 1130 333 1132 335
rect 1096 309 1100 318
rect 1128 317 1132 333
rect 1128 315 1129 317
rect 1131 315 1132 317
rect 1128 314 1132 315
rect 1127 312 1132 314
rect 1127 310 1128 312
rect 1130 310 1132 312
rect 1127 308 1132 310
rect 1087 307 1088 308
rect 1086 306 1088 307
rect 1090 306 1091 308
rect 1086 305 1091 306
rect 1086 303 1087 305
rect 1089 303 1091 305
rect 1086 301 1091 303
rect -290 295 1136 296
rect -290 293 -280 295
rect -278 293 -227 295
rect -225 293 -5 295
rect -3 293 28 295
rect 30 293 38 295
rect 40 293 68 295
rect 70 293 78 295
rect 80 293 297 295
rect 299 293 335 295
rect 337 293 345 295
rect 347 293 574 295
rect 576 293 612 295
rect 614 293 622 295
rect 624 293 850 295
rect 852 293 888 295
rect 890 293 898 295
rect 900 293 1127 295
rect 1129 293 1136 295
rect -290 292 1136 293
rect -290 290 211 292
rect 213 290 488 292
rect 490 290 764 292
rect 766 290 1041 292
rect 1043 290 1136 292
rect -290 288 164 290
rect 166 288 1136 290
rect -287 283 1136 288
rect -287 281 -280 283
rect -278 281 -227 283
rect -225 281 -5 283
rect -3 281 28 283
rect 30 281 38 283
rect 40 281 68 283
rect 70 281 78 283
rect 80 281 297 283
rect 299 281 335 283
rect 337 281 345 283
rect 347 281 574 283
rect 576 281 612 283
rect 614 281 622 283
rect 624 281 850 283
rect 852 281 888 283
rect 890 281 898 283
rect 900 281 1127 283
rect 1129 281 1136 283
rect -287 280 1136 281
rect -247 273 -223 274
rect -247 271 -245 273
rect -243 271 -223 273
rect -247 270 -223 271
rect -275 266 -262 267
rect -275 264 -265 266
rect -263 264 -262 266
rect -275 262 -262 264
rect -275 261 -265 262
rect -267 260 -265 261
rect -263 260 -262 262
rect -283 249 -278 251
rect -283 247 -281 249
rect -279 247 -278 249
rect -283 239 -278 247
rect -267 253 -262 260
rect -227 256 -223 270
rect -227 254 -226 256
rect -224 254 -223 256
rect -283 237 -281 239
rect -279 237 -278 239
rect -283 235 -278 237
rect -283 234 -271 235
rect -288 229 -271 234
rect -227 242 -223 254
rect -239 240 -223 242
rect -239 238 -237 240
rect -235 238 -223 240
rect -239 237 -223 238
rect -215 273 -210 275
rect -215 271 -213 273
rect -211 271 -210 273
rect -215 269 -210 271
rect -215 265 -211 269
rect -215 263 -214 265
rect -212 263 -211 265
rect -215 247 -211 263
rect -136 273 -130 274
rect -136 271 -135 273
rect -133 271 -130 273
rect -136 270 -130 271
rect -215 245 -210 247
rect -215 243 -213 245
rect -211 243 -210 245
rect -215 238 -210 243
rect -187 257 -179 259
rect -167 258 -163 267
rect -187 255 -186 257
rect -184 256 -179 257
rect -184 255 -182 256
rect -187 254 -182 255
rect -180 254 -179 256
rect -169 257 -154 258
rect -169 255 -167 257
rect -165 255 -164 257
rect -162 255 -160 257
rect -158 255 -154 257
rect -169 254 -154 255
rect -187 253 -179 254
rect -184 250 -179 253
rect -134 257 -130 270
rect -134 255 -133 257
rect -131 255 -130 257
rect -184 246 -146 250
rect -134 250 -130 255
rect -136 248 -130 250
rect -136 246 -135 248
rect -133 246 -130 248
rect -136 241 -130 246
rect -136 239 -135 241
rect -133 239 -130 241
rect -215 236 -213 238
rect -211 236 -210 238
rect -215 234 -210 236
rect -136 237 -130 239
rect -126 273 -120 274
rect -126 271 -123 273
rect -121 271 -120 273
rect -126 270 -120 271
rect -46 273 -41 275
rect -46 271 -45 273
rect -43 271 -41 273
rect -126 250 -122 270
rect -93 265 -89 267
rect -93 263 -92 265
rect -90 263 -89 265
rect -126 248 -120 250
rect -126 246 -123 248
rect -121 246 -120 248
rect -126 244 -120 246
rect -126 242 -123 244
rect -121 242 -120 244
rect -126 241 -120 242
rect -126 239 -123 241
rect -121 239 -120 241
rect -126 237 -120 239
rect -93 258 -89 263
rect -46 269 -41 271
rect -45 265 -41 269
rect -45 263 -44 265
rect -42 263 -41 265
rect -102 257 -87 258
rect -102 255 -98 257
rect -96 255 -91 257
rect -89 255 -87 257
rect -102 254 -87 255
rect -77 257 -69 259
rect -77 255 -72 257
rect -70 255 -69 257
rect -77 253 -69 255
rect -77 250 -72 253
rect -110 249 -72 250
rect -110 247 -88 249
rect -86 247 -72 249
rect -110 246 -72 247
rect -45 247 -41 263
rect -36 258 -32 267
rect -36 257 -15 258
rect -36 255 -35 257
rect -33 255 -21 257
rect -19 255 -15 257
rect -36 254 -15 255
rect -5 266 0 268
rect -5 264 -4 266
rect -2 264 0 266
rect -5 262 0 264
rect -46 245 -41 247
rect -46 243 -45 245
rect -43 243 -41 245
rect -46 238 -41 243
rect -46 236 -45 238
rect -43 236 -41 238
rect -36 248 -31 250
rect -29 248 -15 250
rect -36 246 -15 248
rect -36 244 -32 246
rect -36 242 -35 244
rect -33 242 -32 244
rect -4 249 0 262
rect 14 261 19 267
rect 31 271 43 275
rect 31 269 39 271
rect 41 269 43 271
rect 14 259 16 261
rect 18 259 19 261
rect 14 258 19 259
rect 14 257 28 258
rect 14 255 22 257
rect 24 255 28 257
rect 14 254 28 255
rect -4 247 -3 249
rect -1 247 0 249
rect -36 237 -32 242
rect -46 234 -41 236
rect -4 243 0 247
rect -2 241 0 243
rect -4 236 0 241
rect 7 249 20 250
rect 7 247 12 249
rect 14 247 16 249
rect 18 247 20 249
rect 7 246 20 247
rect 7 237 11 246
rect 39 249 43 269
rect 54 266 59 267
rect 54 264 56 266
rect 58 264 59 266
rect 54 258 59 264
rect 71 271 83 275
rect 71 269 79 271
rect 81 269 83 271
rect 54 257 68 258
rect 54 255 62 257
rect 64 255 68 257
rect 54 254 68 255
rect 38 247 40 249
rect 42 247 43 249
rect 38 246 43 247
rect 38 244 39 246
rect 41 244 43 246
rect -2 234 0 236
rect -13 230 0 234
rect -4 229 0 230
rect 38 238 43 244
rect 38 236 39 238
rect 41 236 43 238
rect 47 249 60 250
rect 47 247 52 249
rect 54 247 60 249
rect 47 246 60 247
rect 47 241 51 246
rect 79 257 83 269
rect 79 255 80 257
rect 82 255 83 257
rect 79 249 83 255
rect 47 239 48 241
rect 50 239 51 241
rect 47 237 51 239
rect 78 247 83 249
rect 78 245 79 247
rect 81 245 83 247
rect 78 240 83 245
rect 38 234 43 236
rect 78 238 79 240
rect 81 238 83 240
rect 78 236 83 238
rect 87 273 92 275
rect 87 271 89 273
rect 91 271 92 273
rect 87 269 92 271
rect 87 265 91 269
rect 87 263 88 265
rect 90 263 91 265
rect 87 247 91 263
rect 166 273 172 274
rect 166 271 167 273
rect 169 271 172 273
rect 166 270 172 271
rect 87 245 92 247
rect 87 243 89 245
rect 91 243 92 245
rect 87 238 92 243
rect 115 257 123 259
rect 135 258 139 267
rect 115 255 116 257
rect 118 255 123 257
rect 115 253 123 255
rect 133 257 148 258
rect 133 255 135 257
rect 137 255 138 257
rect 140 255 142 257
rect 144 255 148 257
rect 133 254 148 255
rect 118 250 123 253
rect 168 257 172 270
rect 168 255 169 257
rect 171 255 172 257
rect 118 249 156 250
rect 118 247 133 249
rect 135 247 156 249
rect 118 246 156 247
rect 168 250 172 255
rect 166 248 172 250
rect 166 246 167 248
rect 169 246 172 248
rect 166 241 172 246
rect 166 239 167 241
rect 169 239 172 241
rect 87 236 89 238
rect 91 236 92 238
rect 87 234 92 236
rect 166 237 172 239
rect 176 273 182 274
rect 176 271 179 273
rect 181 271 182 273
rect 176 270 182 271
rect 256 273 263 275
rect 256 271 257 273
rect 259 271 263 273
rect 176 250 180 270
rect 209 265 213 267
rect 209 263 210 265
rect 212 263 213 265
rect 176 248 182 250
rect 176 246 179 248
rect 181 246 182 248
rect 176 244 182 246
rect 176 242 179 244
rect 181 242 182 244
rect 176 241 182 242
rect 176 239 179 241
rect 181 239 182 241
rect 176 237 182 239
rect 209 258 213 263
rect 256 269 260 271
rect 262 269 263 271
rect 257 268 263 269
rect 200 257 215 258
rect 200 255 204 257
rect 206 255 211 257
rect 213 255 215 257
rect 200 254 215 255
rect 225 257 233 259
rect 225 255 230 257
rect 232 255 233 257
rect 225 253 233 255
rect 225 252 230 253
rect 225 250 227 252
rect 229 250 230 252
rect 192 246 230 250
rect 257 247 261 268
rect 266 263 270 264
rect 266 261 267 263
rect 269 261 270 263
rect 266 258 270 261
rect 266 257 287 258
rect 266 255 281 257
rect 283 255 287 257
rect 266 254 287 255
rect 297 266 302 268
rect 297 264 298 266
rect 300 264 302 266
rect 297 262 302 264
rect 256 245 261 247
rect 256 243 257 245
rect 259 243 261 245
rect 256 238 261 243
rect 256 236 257 238
rect 259 236 261 238
rect 266 248 271 250
rect 273 248 287 250
rect 266 246 287 248
rect 266 244 270 246
rect 266 242 267 244
rect 269 242 270 244
rect 266 237 270 242
rect 256 234 261 236
rect 298 243 302 262
rect 321 258 326 267
rect 338 271 350 275
rect 338 269 346 271
rect 348 269 350 271
rect 321 257 335 258
rect 321 255 329 257
rect 331 255 332 257
rect 334 255 335 257
rect 321 254 335 255
rect 300 241 302 243
rect 298 236 302 241
rect 314 249 327 250
rect 314 247 315 249
rect 317 247 319 249
rect 321 247 327 249
rect 314 246 327 247
rect 314 237 318 246
rect 346 256 350 269
rect 346 254 347 256
rect 349 254 350 256
rect 346 249 350 254
rect 345 247 350 249
rect 345 245 346 247
rect 348 245 350 247
rect 345 240 350 245
rect 300 234 302 236
rect 289 233 302 234
rect 289 231 291 233
rect 293 231 302 233
rect 289 230 302 231
rect 298 229 302 230
rect 345 238 346 240
rect 348 238 350 240
rect 345 236 350 238
rect 364 273 369 275
rect 364 271 366 273
rect 368 271 369 273
rect 364 269 369 271
rect 364 265 368 269
rect 364 263 365 265
rect 367 263 368 265
rect 364 247 368 263
rect 443 273 449 274
rect 443 271 444 273
rect 446 271 449 273
rect 443 270 449 271
rect 364 245 369 247
rect 364 243 366 245
rect 368 243 369 245
rect 364 238 369 243
rect 392 257 400 259
rect 412 258 416 267
rect 392 255 393 257
rect 395 255 400 257
rect 392 253 400 255
rect 410 257 425 258
rect 410 255 412 257
rect 414 255 415 257
rect 417 255 419 257
rect 421 255 425 257
rect 410 254 425 255
rect 395 250 400 253
rect 445 257 449 270
rect 445 255 446 257
rect 448 255 449 257
rect 395 249 433 250
rect 395 247 410 249
rect 412 247 433 249
rect 395 246 433 247
rect 445 250 449 255
rect 443 248 449 250
rect 443 246 444 248
rect 446 246 449 248
rect 443 241 449 246
rect 443 239 444 241
rect 446 239 449 241
rect 364 236 366 238
rect 368 236 369 238
rect 364 234 369 236
rect 443 237 449 239
rect 453 273 459 274
rect 453 271 456 273
rect 458 271 459 273
rect 453 270 459 271
rect 533 273 540 275
rect 533 271 534 273
rect 536 271 540 273
rect 453 250 457 270
rect 486 265 490 267
rect 486 263 487 265
rect 489 263 490 265
rect 453 248 459 250
rect 453 246 456 248
rect 458 246 459 248
rect 453 244 459 246
rect 453 242 456 244
rect 458 242 459 244
rect 453 241 459 242
rect 453 239 456 241
rect 458 239 459 241
rect 453 237 459 239
rect 486 258 490 263
rect 533 269 537 271
rect 539 269 540 271
rect 534 268 540 269
rect 477 257 492 258
rect 477 255 481 257
rect 483 255 488 257
rect 490 255 492 257
rect 477 254 492 255
rect 502 257 510 259
rect 502 255 507 257
rect 509 255 510 257
rect 502 253 510 255
rect 502 252 507 253
rect 502 250 504 252
rect 506 250 507 252
rect 469 246 507 250
rect 534 247 538 268
rect 543 263 547 264
rect 543 261 544 263
rect 546 261 547 263
rect 543 258 547 261
rect 543 257 564 258
rect 543 255 558 257
rect 560 255 564 257
rect 543 254 564 255
rect 574 266 579 268
rect 574 264 575 266
rect 577 264 579 266
rect 574 262 579 264
rect 533 245 538 247
rect 533 243 534 245
rect 536 243 538 245
rect 533 238 538 243
rect 533 236 534 238
rect 536 236 538 238
rect 543 248 548 250
rect 550 248 564 250
rect 543 246 564 248
rect 543 244 547 246
rect 543 242 544 244
rect 546 242 547 244
rect 543 237 547 242
rect 533 234 538 236
rect 575 243 579 262
rect 598 258 603 267
rect 615 271 627 275
rect 615 269 623 271
rect 625 269 627 271
rect 598 257 612 258
rect 598 255 606 257
rect 608 255 609 257
rect 611 255 612 257
rect 598 254 612 255
rect 577 241 579 243
rect 575 236 579 241
rect 591 249 604 250
rect 591 247 592 249
rect 594 247 596 249
rect 598 247 604 249
rect 591 246 604 247
rect 591 237 595 246
rect 623 256 627 269
rect 623 254 624 256
rect 626 254 627 256
rect 623 249 627 254
rect 622 247 627 249
rect 622 245 623 247
rect 625 245 627 247
rect 622 240 627 245
rect 577 234 579 236
rect 566 233 579 234
rect 566 231 568 233
rect 570 231 579 233
rect 566 230 579 231
rect 575 229 579 230
rect 622 238 623 240
rect 625 238 627 240
rect 622 236 627 238
rect 640 273 645 275
rect 640 271 642 273
rect 644 271 645 273
rect 640 269 645 271
rect 640 265 644 269
rect 640 263 641 265
rect 643 263 644 265
rect 640 247 644 263
rect 719 273 725 274
rect 719 271 720 273
rect 722 271 725 273
rect 719 270 725 271
rect 640 245 645 247
rect 640 243 642 245
rect 644 243 645 245
rect 640 238 645 243
rect 668 257 676 259
rect 688 258 692 267
rect 668 255 669 257
rect 671 255 676 257
rect 668 253 676 255
rect 686 257 701 258
rect 686 255 688 257
rect 690 255 691 257
rect 693 255 695 257
rect 697 255 701 257
rect 686 254 701 255
rect 671 250 676 253
rect 721 257 725 270
rect 721 255 722 257
rect 724 255 725 257
rect 671 249 709 250
rect 671 247 686 249
rect 688 247 709 249
rect 671 246 709 247
rect 721 250 725 255
rect 719 248 725 250
rect 719 246 720 248
rect 722 246 725 248
rect 719 241 725 246
rect 719 239 720 241
rect 722 239 725 241
rect 640 236 642 238
rect 644 236 645 238
rect 640 234 645 236
rect 719 237 725 239
rect 729 273 735 274
rect 729 271 732 273
rect 734 271 735 273
rect 729 270 735 271
rect 809 273 816 275
rect 809 271 810 273
rect 812 271 816 273
rect 729 250 733 270
rect 762 265 766 267
rect 762 263 763 265
rect 765 263 766 265
rect 729 248 735 250
rect 729 246 732 248
rect 734 246 735 248
rect 729 244 735 246
rect 729 242 732 244
rect 734 242 735 244
rect 729 241 735 242
rect 729 239 732 241
rect 734 239 735 241
rect 729 237 735 239
rect 762 258 766 263
rect 809 269 813 271
rect 815 269 816 271
rect 810 268 816 269
rect 753 257 768 258
rect 753 255 757 257
rect 759 255 764 257
rect 766 255 768 257
rect 753 254 768 255
rect 778 257 786 259
rect 778 255 783 257
rect 785 255 786 257
rect 778 253 786 255
rect 778 252 783 253
rect 778 250 780 252
rect 782 250 783 252
rect 745 246 783 250
rect 810 247 814 268
rect 819 263 823 264
rect 819 261 820 263
rect 822 261 823 263
rect 819 258 823 261
rect 819 257 840 258
rect 819 255 834 257
rect 836 255 840 257
rect 819 254 840 255
rect 850 266 855 268
rect 850 264 851 266
rect 853 264 855 266
rect 850 262 855 264
rect 809 245 814 247
rect 809 243 810 245
rect 812 243 814 245
rect 809 238 814 243
rect 809 236 810 238
rect 812 236 814 238
rect 819 248 824 250
rect 826 248 840 250
rect 819 246 840 248
rect 819 244 823 246
rect 819 242 820 244
rect 822 242 823 244
rect 819 237 823 242
rect 809 234 814 236
rect 851 243 855 262
rect 874 258 879 267
rect 891 271 903 275
rect 891 269 899 271
rect 901 269 903 271
rect 874 257 888 258
rect 874 255 882 257
rect 884 255 885 257
rect 887 255 888 257
rect 874 254 888 255
rect 853 241 855 243
rect 851 236 855 241
rect 867 249 880 250
rect 867 247 868 249
rect 870 247 872 249
rect 874 247 880 249
rect 867 246 880 247
rect 867 237 871 246
rect 899 256 903 269
rect 899 254 900 256
rect 902 254 903 256
rect 899 249 903 254
rect 898 247 903 249
rect 898 245 899 247
rect 901 245 903 247
rect 898 240 903 245
rect 853 234 855 236
rect 842 233 855 234
rect 842 231 844 233
rect 846 231 855 233
rect 842 230 855 231
rect 851 229 855 230
rect 898 238 899 240
rect 901 238 903 240
rect 898 236 903 238
rect 917 273 922 275
rect 917 271 919 273
rect 921 271 922 273
rect 917 269 922 271
rect 917 265 921 269
rect 917 263 918 265
rect 920 263 921 265
rect 917 247 921 263
rect 996 273 1002 274
rect 996 271 997 273
rect 999 271 1002 273
rect 996 270 1002 271
rect 917 245 922 247
rect 917 243 919 245
rect 921 243 922 245
rect 917 238 922 243
rect 945 257 953 259
rect 965 258 969 267
rect 945 255 946 257
rect 948 255 953 257
rect 945 253 953 255
rect 963 257 978 258
rect 963 255 965 257
rect 967 255 968 257
rect 970 255 972 257
rect 974 255 978 257
rect 963 254 978 255
rect 948 250 953 253
rect 998 257 1002 270
rect 998 255 999 257
rect 1001 255 1002 257
rect 948 249 986 250
rect 948 247 963 249
rect 965 247 986 249
rect 948 246 986 247
rect 998 250 1002 255
rect 996 248 1002 250
rect 996 246 997 248
rect 999 246 1002 248
rect 996 241 1002 246
rect 996 239 997 241
rect 999 239 1002 241
rect 917 236 919 238
rect 921 236 922 238
rect 917 234 922 236
rect 996 237 1002 239
rect 1006 273 1012 274
rect 1006 271 1009 273
rect 1011 271 1012 273
rect 1006 270 1012 271
rect 1086 274 1093 275
rect 1086 273 1090 274
rect 1086 271 1087 273
rect 1089 272 1090 273
rect 1092 272 1093 274
rect 1089 271 1093 272
rect 1006 250 1010 270
rect 1039 265 1043 267
rect 1039 263 1040 265
rect 1042 263 1043 265
rect 1006 248 1012 250
rect 1006 246 1009 248
rect 1011 246 1012 248
rect 1006 244 1012 246
rect 1006 242 1009 244
rect 1011 242 1012 244
rect 1006 241 1012 242
rect 1006 239 1009 241
rect 1011 239 1012 241
rect 1006 237 1012 239
rect 1039 258 1043 263
rect 1086 269 1093 271
rect 1087 268 1093 269
rect 1030 257 1045 258
rect 1030 255 1034 257
rect 1036 255 1041 257
rect 1043 255 1045 257
rect 1030 254 1045 255
rect 1055 257 1063 259
rect 1055 255 1060 257
rect 1062 255 1063 257
rect 1055 253 1063 255
rect 1055 252 1060 253
rect 1055 250 1057 252
rect 1059 250 1060 252
rect 1022 246 1060 250
rect 1087 247 1091 268
rect 1096 263 1100 264
rect 1096 261 1097 263
rect 1099 261 1100 263
rect 1096 258 1100 261
rect 1096 257 1117 258
rect 1096 255 1111 257
rect 1113 255 1117 257
rect 1096 254 1117 255
rect 1127 266 1132 268
rect 1127 264 1128 266
rect 1130 264 1132 266
rect 1127 262 1132 264
rect 1086 245 1091 247
rect 1086 243 1087 245
rect 1089 243 1091 245
rect 1086 238 1091 243
rect 1086 236 1087 238
rect 1089 236 1091 238
rect 1096 248 1101 250
rect 1103 248 1117 250
rect 1096 246 1117 248
rect 1096 244 1100 246
rect 1096 242 1097 244
rect 1099 242 1100 244
rect 1096 237 1100 242
rect 1086 234 1091 236
rect 1128 243 1132 262
rect 1130 241 1132 243
rect 1128 236 1132 241
rect 1130 234 1132 236
rect 1119 233 1132 234
rect 1119 231 1121 233
rect 1123 231 1132 233
rect 1119 230 1132 231
rect 1128 229 1132 230
rect -287 223 1136 224
rect -287 221 -247 223
rect -245 221 -5 223
rect -3 221 38 223
rect 40 221 78 223
rect 80 221 297 223
rect 299 221 345 223
rect 347 221 574 223
rect 576 221 622 223
rect 624 221 850 223
rect 852 221 898 223
rect 900 221 1127 223
rect 1129 221 1136 223
rect -287 218 1136 221
rect -287 216 100 218
rect 102 216 1136 218
rect -287 211 1136 216
rect -287 209 -247 211
rect -245 209 -5 211
rect -3 209 38 211
rect 40 209 78 211
rect 80 209 297 211
rect 299 209 345 211
rect 347 209 574 211
rect 576 209 622 211
rect 624 209 850 211
rect 852 209 898 211
rect 900 209 1127 211
rect 1129 209 1136 211
rect -287 208 1136 209
rect -283 197 -271 203
rect -283 196 -278 197
rect -286 189 -278 196
rect -283 188 -278 189
rect -4 202 0 203
rect -13 198 0 202
rect -215 196 -210 198
rect -283 186 -281 188
rect -279 186 -278 188
rect -283 185 -278 186
rect -283 183 -281 185
rect -279 183 -278 185
rect -283 181 -278 183
rect -267 177 -262 179
rect -267 175 -265 177
rect -263 175 -262 177
rect -267 172 -262 175
rect -239 194 -223 195
rect -239 192 -237 194
rect -235 192 -223 194
rect -239 190 -223 192
rect -227 178 -223 190
rect -227 176 -226 178
rect -224 176 -223 178
rect -267 171 -265 172
rect -275 170 -265 171
rect -263 170 -262 172
rect -275 165 -262 170
rect -227 162 -223 176
rect -247 161 -223 162
rect -247 159 -245 161
rect -243 159 -223 161
rect -247 158 -223 159
rect -215 194 -213 196
rect -211 194 -210 196
rect -215 189 -210 194
rect -215 187 -213 189
rect -211 187 -210 189
rect -215 185 -210 187
rect -215 169 -211 185
rect -184 182 -146 186
rect -184 179 -179 182
rect -187 178 -179 179
rect -187 177 -182 178
rect -187 175 -186 177
rect -184 176 -182 177
rect -180 176 -179 178
rect -184 175 -179 176
rect -187 173 -179 175
rect -169 177 -154 178
rect -169 175 -167 177
rect -165 175 -163 177
rect -161 175 -160 177
rect -158 175 -154 177
rect -169 174 -154 175
rect -215 167 -214 169
rect -212 167 -211 169
rect -215 163 -211 167
rect -215 161 -210 163
rect -167 165 -163 174
rect -136 193 -130 195
rect -136 191 -135 193
rect -133 191 -130 193
rect -136 186 -130 191
rect -136 184 -135 186
rect -133 184 -130 186
rect -136 182 -130 184
rect -134 177 -130 182
rect -134 175 -133 177
rect -131 175 -130 177
rect -134 162 -130 175
rect -215 159 -213 161
rect -211 159 -210 161
rect -215 157 -210 159
rect -136 161 -130 162
rect -136 159 -135 161
rect -133 159 -130 161
rect -136 158 -130 159
rect -126 193 -120 195
rect -46 196 -41 198
rect -46 194 -45 196
rect -43 194 -41 196
rect -126 191 -123 193
rect -121 191 -120 193
rect -126 190 -120 191
rect -126 188 -123 190
rect -121 188 -120 190
rect -126 186 -120 188
rect -126 184 -123 186
rect -121 184 -120 186
rect -126 182 -120 184
rect -126 162 -122 182
rect -110 185 -72 186
rect -110 183 -86 185
rect -84 183 -72 185
rect -110 182 -72 183
rect -77 179 -72 182
rect -102 177 -87 178
rect -102 175 -98 177
rect -96 175 -91 177
rect -89 175 -87 177
rect -102 174 -87 175
rect -77 177 -69 179
rect -77 175 -72 177
rect -70 175 -69 177
rect -93 169 -89 174
rect -77 173 -69 175
rect -46 189 -41 194
rect -46 187 -45 189
rect -43 187 -41 189
rect -46 185 -41 187
rect -93 167 -92 169
rect -90 167 -89 169
rect -93 165 -89 167
rect -126 161 -120 162
rect -126 159 -123 161
rect -121 159 -120 161
rect -126 158 -120 159
rect -45 167 -41 185
rect -36 190 -32 195
rect -36 188 -35 190
rect -33 188 -32 190
rect -36 186 -32 188
rect -36 184 -15 186
rect -36 182 -31 184
rect -29 182 -15 184
rect -45 165 -44 167
rect -42 165 -41 167
rect -36 177 -15 178
rect -36 175 -35 177
rect -33 175 -21 177
rect -19 175 -15 177
rect -36 174 -15 175
rect -2 196 0 198
rect -4 191 0 196
rect -2 189 0 191
rect -36 165 -32 174
rect -4 173 0 189
rect 7 188 11 195
rect 38 197 43 199
rect 38 195 39 197
rect 41 195 43 197
rect 7 186 8 188
rect 10 186 11 188
rect 7 185 20 186
rect 7 183 12 185
rect 14 183 20 185
rect 7 182 20 183
rect -4 171 -3 173
rect -1 171 0 173
rect -4 170 0 171
rect -5 168 0 170
rect -5 166 -4 168
rect -2 166 0 168
rect -45 163 -41 165
rect -5 164 0 166
rect 14 177 28 178
rect 14 175 22 177
rect 24 175 28 177
rect 14 174 28 175
rect 38 189 43 195
rect 38 187 39 189
rect 41 187 43 189
rect 38 185 43 187
rect 38 183 40 185
rect 42 183 43 185
rect 38 181 43 183
rect 47 194 51 195
rect 47 192 48 194
rect 50 192 51 194
rect 47 186 51 192
rect 298 202 302 203
rect 289 198 302 202
rect 87 196 92 198
rect 78 194 83 196
rect 47 185 60 186
rect 47 183 52 185
rect 54 183 60 185
rect 47 182 60 183
rect 14 169 19 174
rect 14 167 16 169
rect 18 167 19 169
rect 14 165 19 167
rect -46 161 -41 163
rect 39 163 43 181
rect 54 177 68 178
rect 54 175 62 177
rect 64 175 68 177
rect 54 174 68 175
rect 78 192 79 194
rect 81 192 83 194
rect 78 187 83 192
rect 78 185 79 187
rect 81 185 83 187
rect 78 183 83 185
rect 54 172 59 174
rect 54 170 56 172
rect 58 170 59 172
rect 54 165 59 170
rect 79 177 83 183
rect 79 175 80 177
rect 82 175 83 177
rect -46 159 -45 161
rect -43 159 -41 161
rect -46 157 -41 159
rect 31 161 39 163
rect 41 161 43 163
rect 79 163 83 175
rect 31 157 43 161
rect 71 161 79 163
rect 81 161 83 163
rect 71 157 83 161
rect 87 194 89 196
rect 91 194 92 196
rect 87 189 92 194
rect 87 187 89 189
rect 91 187 92 189
rect 87 185 92 187
rect 87 169 91 185
rect 118 185 156 186
rect 118 183 137 185
rect 139 183 156 185
rect 118 182 156 183
rect 118 179 123 182
rect 115 177 123 179
rect 115 175 116 177
rect 118 175 123 177
rect 115 173 123 175
rect 133 177 148 178
rect 133 175 135 177
rect 137 175 139 177
rect 141 175 142 177
rect 144 175 148 177
rect 133 174 148 175
rect 87 167 88 169
rect 90 167 91 169
rect 87 163 91 167
rect 87 161 92 163
rect 135 165 139 174
rect 166 193 172 195
rect 166 191 167 193
rect 169 191 172 193
rect 166 186 172 191
rect 166 184 167 186
rect 169 184 172 186
rect 166 182 172 184
rect 168 177 172 182
rect 168 175 169 177
rect 171 175 172 177
rect 168 162 172 175
rect 87 159 89 161
rect 91 159 92 161
rect 87 157 92 159
rect 166 161 172 162
rect 166 159 167 161
rect 169 159 172 161
rect 166 158 172 159
rect 176 193 182 195
rect 256 196 261 198
rect 256 194 257 196
rect 259 194 261 196
rect 176 191 179 193
rect 181 191 182 193
rect 176 190 182 191
rect 176 188 179 190
rect 181 188 182 190
rect 176 186 182 188
rect 176 184 179 186
rect 181 184 182 186
rect 176 182 182 184
rect 176 162 180 182
rect 192 185 230 186
rect 192 183 227 185
rect 229 183 230 185
rect 192 182 230 183
rect 225 179 230 182
rect 200 177 215 178
rect 200 175 204 177
rect 206 175 211 177
rect 213 175 215 177
rect 200 174 215 175
rect 225 177 233 179
rect 225 175 230 177
rect 232 175 233 177
rect 209 169 213 174
rect 225 173 233 175
rect 256 189 261 194
rect 256 187 257 189
rect 259 187 261 189
rect 256 185 261 187
rect 209 167 210 169
rect 212 167 213 169
rect 209 165 213 167
rect 176 161 182 162
rect 176 159 179 161
rect 181 159 182 161
rect 176 158 182 159
rect 257 163 261 185
rect 266 194 270 195
rect 266 192 267 194
rect 269 192 270 194
rect 266 186 270 192
rect 266 184 287 186
rect 266 182 271 184
rect 273 182 287 184
rect 266 177 287 178
rect 266 175 267 177
rect 269 175 281 177
rect 283 175 287 177
rect 266 174 287 175
rect 300 196 302 198
rect 298 191 302 196
rect 300 189 302 191
rect 266 170 270 174
rect 298 173 302 189
rect 314 189 318 195
rect 575 202 579 203
rect 566 198 579 202
rect 364 196 369 198
rect 345 194 350 196
rect 314 187 315 189
rect 317 187 318 189
rect 314 186 318 187
rect 314 185 327 186
rect 314 183 319 185
rect 321 183 327 185
rect 314 182 327 183
rect 298 171 299 173
rect 301 171 302 173
rect 298 170 302 171
rect 297 168 302 170
rect 297 166 298 168
rect 300 166 302 168
rect 297 164 302 166
rect 321 177 335 178
rect 321 175 329 177
rect 331 175 332 177
rect 334 175 335 177
rect 321 174 335 175
rect 345 192 346 194
rect 348 192 350 194
rect 345 187 350 192
rect 345 185 346 187
rect 348 185 350 187
rect 345 183 350 185
rect 321 165 326 174
rect 346 182 350 183
rect 346 180 347 182
rect 349 180 350 182
rect 256 161 263 163
rect 346 163 350 180
rect 256 159 257 161
rect 259 159 260 161
rect 262 159 263 161
rect 256 157 263 159
rect 338 161 346 163
rect 348 161 350 163
rect 338 157 350 161
rect 364 194 366 196
rect 368 194 369 196
rect 364 189 369 194
rect 364 187 366 189
rect 368 187 369 189
rect 364 185 369 187
rect 364 169 368 185
rect 395 185 433 186
rect 395 183 414 185
rect 416 183 433 185
rect 395 182 433 183
rect 395 179 400 182
rect 392 177 400 179
rect 392 175 393 177
rect 395 175 400 177
rect 392 173 400 175
rect 410 177 425 178
rect 410 175 412 177
rect 414 175 416 177
rect 418 175 419 177
rect 421 175 425 177
rect 410 174 425 175
rect 364 167 365 169
rect 367 167 368 169
rect 364 163 368 167
rect 364 161 369 163
rect 412 165 416 174
rect 443 193 449 195
rect 443 191 444 193
rect 446 191 449 193
rect 443 186 449 191
rect 443 184 444 186
rect 446 184 449 186
rect 443 182 449 184
rect 445 177 449 182
rect 445 175 446 177
rect 448 175 449 177
rect 445 162 449 175
rect 364 159 366 161
rect 368 159 369 161
rect 364 157 369 159
rect 443 161 449 162
rect 443 159 444 161
rect 446 159 449 161
rect 443 158 449 159
rect 453 193 459 195
rect 533 196 538 198
rect 533 194 534 196
rect 536 194 538 196
rect 453 191 456 193
rect 458 191 459 193
rect 453 190 459 191
rect 453 188 456 190
rect 458 188 459 190
rect 453 186 459 188
rect 453 184 456 186
rect 458 184 459 186
rect 453 182 459 184
rect 453 162 457 182
rect 469 185 507 186
rect 469 183 504 185
rect 506 183 507 185
rect 469 182 507 183
rect 502 179 507 182
rect 477 177 492 178
rect 477 175 481 177
rect 483 175 488 177
rect 490 175 492 177
rect 477 174 492 175
rect 502 177 510 179
rect 502 175 507 177
rect 509 175 510 177
rect 486 169 490 174
rect 502 173 510 175
rect 533 189 538 194
rect 533 187 534 189
rect 536 187 538 189
rect 533 185 538 187
rect 486 167 487 169
rect 489 167 490 169
rect 486 165 490 167
rect 453 161 459 162
rect 453 159 456 161
rect 458 159 459 161
rect 453 158 459 159
rect 534 163 538 185
rect 543 194 547 195
rect 543 192 544 194
rect 546 192 547 194
rect 543 186 547 192
rect 543 184 564 186
rect 543 182 548 184
rect 550 182 564 184
rect 543 177 564 178
rect 543 175 544 177
rect 546 175 558 177
rect 560 175 564 177
rect 543 174 564 175
rect 577 196 579 198
rect 575 191 579 196
rect 577 189 579 191
rect 543 170 547 174
rect 575 173 579 189
rect 591 189 595 195
rect 851 202 855 203
rect 842 198 855 202
rect 640 196 645 198
rect 622 194 627 196
rect 591 187 592 189
rect 594 187 595 189
rect 591 186 595 187
rect 591 185 604 186
rect 591 183 596 185
rect 598 183 604 185
rect 591 182 604 183
rect 575 171 576 173
rect 578 171 579 173
rect 575 170 579 171
rect 574 168 579 170
rect 574 166 575 168
rect 577 166 579 168
rect 574 164 579 166
rect 598 177 612 178
rect 598 175 606 177
rect 608 175 609 177
rect 611 175 612 177
rect 598 174 612 175
rect 622 192 623 194
rect 625 192 627 194
rect 622 187 627 192
rect 622 185 623 187
rect 625 185 627 187
rect 622 183 627 185
rect 598 165 603 174
rect 623 182 627 183
rect 623 180 624 182
rect 626 180 627 182
rect 533 161 540 163
rect 623 163 627 180
rect 533 159 534 161
rect 536 159 537 161
rect 539 159 540 161
rect 533 157 540 159
rect 615 161 623 163
rect 625 161 627 163
rect 615 157 627 161
rect 640 194 642 196
rect 644 194 645 196
rect 640 189 645 194
rect 640 187 642 189
rect 644 187 645 189
rect 640 185 645 187
rect 640 169 644 185
rect 671 185 709 186
rect 671 183 690 185
rect 692 183 709 185
rect 671 182 709 183
rect 671 179 676 182
rect 668 177 676 179
rect 668 175 669 177
rect 671 175 676 177
rect 668 173 676 175
rect 686 177 701 178
rect 686 175 688 177
rect 690 175 692 177
rect 694 175 695 177
rect 697 175 701 177
rect 686 174 701 175
rect 640 167 641 169
rect 643 167 644 169
rect 640 163 644 167
rect 640 161 645 163
rect 688 165 692 174
rect 719 193 725 195
rect 719 191 720 193
rect 722 191 725 193
rect 719 186 725 191
rect 719 184 720 186
rect 722 184 725 186
rect 719 182 725 184
rect 721 177 725 182
rect 721 175 722 177
rect 724 175 725 177
rect 721 162 725 175
rect 640 159 642 161
rect 644 159 645 161
rect 640 157 645 159
rect 719 161 725 162
rect 719 159 720 161
rect 722 159 725 161
rect 719 158 725 159
rect 729 193 735 195
rect 809 196 814 198
rect 809 194 810 196
rect 812 194 814 196
rect 729 191 732 193
rect 734 191 735 193
rect 729 190 735 191
rect 729 188 732 190
rect 734 188 735 190
rect 729 186 735 188
rect 729 184 732 186
rect 734 184 735 186
rect 729 182 735 184
rect 729 162 733 182
rect 745 185 783 186
rect 745 183 780 185
rect 782 183 783 185
rect 745 182 783 183
rect 778 179 783 182
rect 753 177 768 178
rect 753 175 757 177
rect 759 175 764 177
rect 766 175 768 177
rect 753 174 768 175
rect 778 177 786 179
rect 778 175 783 177
rect 785 175 786 177
rect 762 169 766 174
rect 778 173 786 175
rect 809 189 814 194
rect 809 187 810 189
rect 812 187 814 189
rect 809 185 814 187
rect 762 167 763 169
rect 765 167 766 169
rect 762 165 766 167
rect 729 161 735 162
rect 729 159 732 161
rect 734 159 735 161
rect 729 158 735 159
rect 810 163 814 185
rect 819 194 823 195
rect 819 192 820 194
rect 822 192 823 194
rect 819 186 823 192
rect 819 184 840 186
rect 819 182 824 184
rect 826 182 840 184
rect 819 177 840 178
rect 819 175 820 177
rect 822 175 834 177
rect 836 175 840 177
rect 819 174 840 175
rect 853 196 855 198
rect 851 191 855 196
rect 853 189 855 191
rect 819 170 823 174
rect 851 173 855 189
rect 867 189 871 195
rect 1128 202 1132 203
rect 1119 198 1132 202
rect 917 196 922 198
rect 898 194 903 196
rect 867 187 868 189
rect 870 187 871 189
rect 867 186 871 187
rect 867 185 880 186
rect 867 183 872 185
rect 874 183 880 185
rect 867 182 880 183
rect 851 171 852 173
rect 854 171 855 173
rect 851 170 855 171
rect 850 168 855 170
rect 850 166 851 168
rect 853 166 855 168
rect 850 164 855 166
rect 874 177 888 178
rect 874 175 882 177
rect 884 175 885 177
rect 887 175 888 177
rect 874 174 888 175
rect 898 192 899 194
rect 901 192 903 194
rect 898 187 903 192
rect 898 185 899 187
rect 901 185 903 187
rect 898 183 903 185
rect 874 165 879 174
rect 899 182 903 183
rect 899 180 900 182
rect 902 180 903 182
rect 809 161 816 163
rect 899 163 903 180
rect 809 159 810 161
rect 812 159 813 161
rect 815 159 816 161
rect 809 157 816 159
rect 891 161 899 163
rect 901 161 903 163
rect 891 157 903 161
rect 917 194 919 196
rect 921 194 922 196
rect 917 189 922 194
rect 917 187 919 189
rect 921 187 922 189
rect 917 185 922 187
rect 917 169 921 185
rect 948 185 986 186
rect 948 183 967 185
rect 969 183 986 185
rect 948 182 986 183
rect 948 179 953 182
rect 945 177 953 179
rect 945 175 946 177
rect 948 175 953 177
rect 945 173 953 175
rect 963 177 978 178
rect 963 175 965 177
rect 967 175 969 177
rect 971 175 972 177
rect 974 175 978 177
rect 963 174 978 175
rect 917 167 918 169
rect 920 167 921 169
rect 917 163 921 167
rect 917 161 922 163
rect 965 165 969 174
rect 996 193 1002 195
rect 996 191 997 193
rect 999 191 1002 193
rect 996 186 1002 191
rect 996 184 997 186
rect 999 184 1002 186
rect 996 182 1002 184
rect 998 177 1002 182
rect 998 175 999 177
rect 1001 175 1002 177
rect 998 162 1002 175
rect 917 159 919 161
rect 921 159 922 161
rect 917 157 922 159
rect 996 161 1002 162
rect 996 159 997 161
rect 999 159 1002 161
rect 996 158 1002 159
rect 1006 193 1012 195
rect 1086 196 1091 198
rect 1086 194 1087 196
rect 1089 194 1091 196
rect 1006 191 1009 193
rect 1011 191 1012 193
rect 1006 190 1012 191
rect 1006 188 1009 190
rect 1011 188 1012 190
rect 1006 186 1012 188
rect 1006 184 1009 186
rect 1011 184 1012 186
rect 1006 182 1012 184
rect 1006 162 1010 182
rect 1022 185 1060 186
rect 1022 183 1057 185
rect 1059 183 1060 185
rect 1022 182 1060 183
rect 1055 179 1060 182
rect 1030 177 1045 178
rect 1030 175 1034 177
rect 1036 175 1041 177
rect 1043 175 1045 177
rect 1030 174 1045 175
rect 1055 177 1063 179
rect 1055 175 1060 177
rect 1062 175 1063 177
rect 1039 169 1043 174
rect 1055 173 1063 175
rect 1086 189 1091 194
rect 1086 187 1087 189
rect 1089 187 1091 189
rect 1086 185 1091 187
rect 1039 167 1040 169
rect 1042 167 1043 169
rect 1039 165 1043 167
rect 1006 161 1012 162
rect 1006 159 1009 161
rect 1011 159 1012 161
rect 1006 158 1012 159
rect 1087 164 1091 185
rect 1096 194 1100 195
rect 1096 192 1097 194
rect 1099 192 1100 194
rect 1096 186 1100 192
rect 1096 184 1117 186
rect 1096 182 1101 184
rect 1103 182 1117 184
rect 1096 177 1117 178
rect 1096 175 1097 177
rect 1099 175 1111 177
rect 1113 175 1117 177
rect 1096 174 1117 175
rect 1130 196 1132 198
rect 1128 191 1132 196
rect 1130 189 1132 191
rect 1096 170 1100 174
rect 1128 173 1132 189
rect 1128 171 1129 173
rect 1131 171 1132 173
rect 1128 170 1132 171
rect 1127 168 1132 170
rect 1127 166 1128 168
rect 1130 166 1132 168
rect 1127 164 1132 166
rect 1087 163 1088 164
rect 1086 162 1088 163
rect 1090 163 1091 164
rect 1090 162 1093 163
rect 1086 161 1093 162
rect 1086 159 1087 161
rect 1089 159 1093 161
rect 1086 157 1093 159
rect -287 151 1136 152
rect -287 149 -280 151
rect -278 149 -227 151
rect -225 149 -5 151
rect -3 149 28 151
rect 30 149 38 151
rect 40 149 68 151
rect 70 149 78 151
rect 80 149 297 151
rect 299 149 335 151
rect 337 149 345 151
rect 347 149 574 151
rect 576 149 612 151
rect 614 149 622 151
rect 624 149 850 151
rect 852 149 888 151
rect 890 149 898 151
rect 900 149 1127 151
rect 1129 149 1136 151
rect -287 146 1136 149
rect -287 144 165 146
rect 167 144 1136 146
rect -287 139 1136 144
rect -287 137 -280 139
rect -278 137 -227 139
rect -225 137 -5 139
rect -3 137 28 139
rect 30 137 38 139
rect 40 137 68 139
rect 70 137 78 139
rect 80 137 297 139
rect 299 137 335 139
rect 337 137 345 139
rect 347 137 574 139
rect 576 137 612 139
rect 614 137 622 139
rect 624 137 850 139
rect 852 137 888 139
rect 890 137 898 139
rect 900 137 1127 139
rect 1129 137 1136 139
rect -287 136 1136 137
rect -247 129 -223 130
rect -247 127 -245 129
rect -243 127 -223 129
rect -247 126 -223 127
rect -275 122 -262 123
rect -275 120 -265 122
rect -263 120 -262 122
rect -275 118 -262 120
rect -275 117 -265 118
rect -267 116 -265 117
rect -263 116 -262 118
rect -283 105 -278 107
rect -283 103 -281 105
rect -279 103 -278 105
rect -283 100 -278 103
rect -267 109 -262 116
rect -227 112 -223 126
rect -227 110 -226 112
rect -224 110 -223 112
rect -289 93 -278 100
rect -283 92 -278 93
rect -283 90 -281 92
rect -279 91 -278 92
rect -279 90 -271 91
rect -283 85 -271 90
rect -227 98 -223 110
rect -239 96 -223 98
rect -239 94 -237 96
rect -235 94 -223 96
rect -239 93 -223 94
rect -215 129 -210 131
rect -215 127 -213 129
rect -211 127 -210 129
rect -215 125 -210 127
rect -215 121 -211 125
rect -215 119 -214 121
rect -212 119 -211 121
rect -215 103 -211 119
rect -136 129 -130 130
rect -136 127 -135 129
rect -133 127 -130 129
rect -136 126 -130 127
rect -215 101 -210 103
rect -215 99 -213 101
rect -211 99 -210 101
rect -215 94 -210 99
rect -187 113 -179 115
rect -167 114 -163 123
rect -187 111 -186 113
rect -184 112 -179 113
rect -184 111 -182 112
rect -187 110 -182 111
rect -180 110 -179 112
rect -169 113 -154 114
rect -169 111 -167 113
rect -165 111 -160 113
rect -158 111 -157 113
rect -155 111 -154 113
rect -169 110 -154 111
rect -187 109 -179 110
rect -184 106 -179 109
rect -134 113 -130 126
rect -134 111 -133 113
rect -131 111 -130 113
rect -184 102 -146 106
rect -134 106 -130 111
rect -136 104 -130 106
rect -136 102 -135 104
rect -133 102 -130 104
rect -136 97 -130 102
rect -136 95 -135 97
rect -133 95 -130 97
rect -215 92 -213 94
rect -211 92 -210 94
rect -215 90 -210 92
rect -136 93 -130 95
rect -126 129 -120 130
rect -126 127 -123 129
rect -121 127 -120 129
rect -126 126 -120 127
rect -46 129 -41 131
rect -46 127 -45 129
rect -43 127 -41 129
rect -126 106 -122 126
rect -93 121 -89 123
rect -93 119 -92 121
rect -90 119 -89 121
rect -126 104 -120 106
rect -126 102 -123 104
rect -121 102 -120 104
rect -126 100 -120 102
rect -126 98 -123 100
rect -121 98 -120 100
rect -126 97 -120 98
rect -126 95 -123 97
rect -121 95 -120 97
rect -126 93 -120 95
rect -93 114 -89 119
rect -46 126 -41 127
rect -46 125 -44 126
rect -45 124 -44 125
rect -42 124 -41 126
rect -102 113 -87 114
rect -102 111 -98 113
rect -96 111 -91 113
rect -89 111 -87 113
rect -102 110 -87 111
rect -77 113 -69 115
rect -77 111 -72 113
rect -70 111 -69 113
rect -77 109 -69 111
rect -77 106 -72 109
rect -110 105 -72 106
rect -110 103 -88 105
rect -86 103 -72 105
rect -110 102 -72 103
rect -45 103 -41 124
rect -36 114 -32 123
rect -36 113 -15 114
rect -36 111 -35 113
rect -33 111 -21 113
rect -19 111 -15 113
rect -36 110 -15 111
rect -5 122 0 124
rect -5 120 -4 122
rect -2 120 0 122
rect -5 118 0 120
rect -46 101 -41 103
rect -46 99 -45 101
rect -43 99 -41 101
rect -46 94 -41 99
rect -46 92 -45 94
rect -43 92 -41 94
rect -36 104 -31 106
rect -29 104 -15 106
rect -36 102 -15 104
rect -36 100 -32 102
rect -36 98 -35 100
rect -33 98 -32 100
rect -4 105 0 118
rect 14 117 19 123
rect 31 127 43 131
rect 31 125 39 127
rect 41 125 43 127
rect 14 115 16 117
rect 18 115 19 117
rect 14 114 19 115
rect 14 113 28 114
rect 14 111 22 113
rect 24 111 28 113
rect 14 110 28 111
rect -4 103 -3 105
rect -1 103 0 105
rect -36 93 -32 98
rect -46 90 -41 92
rect -4 99 0 103
rect -2 97 0 99
rect -4 92 0 97
rect 7 105 20 106
rect 7 103 12 105
rect 14 103 17 105
rect 19 103 20 105
rect 7 102 20 103
rect 7 93 11 102
rect 39 105 43 125
rect 54 121 59 123
rect 54 119 56 121
rect 58 119 59 121
rect 54 114 59 119
rect 71 127 83 131
rect 71 125 79 127
rect 81 125 83 127
rect 54 113 68 114
rect 54 111 62 113
rect 64 111 68 113
rect 54 110 68 111
rect 38 103 40 105
rect 42 103 43 105
rect 38 100 43 103
rect 38 98 39 100
rect 41 98 43 100
rect -2 90 0 92
rect -13 86 0 90
rect -4 85 0 86
rect 38 93 43 98
rect 47 105 60 106
rect 47 103 52 105
rect 54 103 60 105
rect 47 102 60 103
rect 47 97 51 102
rect 79 113 83 125
rect 79 111 80 113
rect 82 111 83 113
rect 79 105 83 111
rect 47 95 48 97
rect 50 95 51 97
rect 47 94 51 95
rect 78 103 83 105
rect 78 101 79 103
rect 81 101 83 103
rect 78 96 83 101
rect 38 91 39 93
rect 41 91 43 93
rect 38 89 43 91
rect 78 94 79 96
rect 81 94 83 96
rect 78 92 83 94
rect 87 129 92 131
rect 87 127 89 129
rect 91 127 92 129
rect 87 125 92 127
rect 87 121 91 125
rect 87 119 88 121
rect 90 119 91 121
rect 87 103 91 119
rect 166 129 172 130
rect 166 127 167 129
rect 169 127 172 129
rect 166 126 172 127
rect 87 101 92 103
rect 87 99 89 101
rect 91 99 92 101
rect 87 94 92 99
rect 115 113 123 115
rect 135 114 139 123
rect 115 111 116 113
rect 118 111 123 113
rect 115 109 123 111
rect 133 113 148 114
rect 133 111 135 113
rect 137 111 138 113
rect 140 111 142 113
rect 144 111 148 113
rect 133 110 148 111
rect 118 106 123 109
rect 168 113 172 126
rect 168 111 169 113
rect 171 111 172 113
rect 118 105 156 106
rect 118 103 131 105
rect 133 103 156 105
rect 118 102 156 103
rect 168 106 172 111
rect 166 104 172 106
rect 166 102 167 104
rect 169 102 172 104
rect 166 97 172 102
rect 166 95 167 97
rect 169 95 172 97
rect 87 92 89 94
rect 91 92 92 94
rect 87 90 92 92
rect 166 93 172 95
rect 176 129 182 130
rect 176 127 179 129
rect 181 127 182 129
rect 176 126 182 127
rect 256 129 263 131
rect 256 127 257 129
rect 259 127 263 129
rect 176 106 180 126
rect 209 121 213 123
rect 209 119 210 121
rect 212 119 213 121
rect 176 104 182 106
rect 176 102 179 104
rect 181 102 182 104
rect 176 100 182 102
rect 176 98 179 100
rect 181 98 182 100
rect 176 97 182 98
rect 176 95 179 97
rect 181 95 182 97
rect 176 93 182 95
rect 209 114 213 119
rect 256 125 260 127
rect 262 125 263 127
rect 257 124 263 125
rect 200 113 215 114
rect 200 111 204 113
rect 206 111 211 113
rect 213 111 215 113
rect 200 110 215 111
rect 225 113 233 115
rect 225 111 230 113
rect 232 111 233 113
rect 225 109 233 111
rect 225 108 230 109
rect 225 106 227 108
rect 229 106 230 108
rect 192 102 230 106
rect 257 103 261 124
rect 266 119 270 120
rect 266 117 267 119
rect 269 117 270 119
rect 266 114 270 117
rect 266 113 287 114
rect 266 111 281 113
rect 283 111 287 113
rect 266 110 287 111
rect 297 122 302 124
rect 297 120 298 122
rect 300 120 302 122
rect 297 118 302 120
rect 256 101 261 103
rect 256 99 257 101
rect 259 99 261 101
rect 256 94 261 99
rect 256 92 257 94
rect 259 92 261 94
rect 266 104 271 106
rect 273 104 287 106
rect 266 102 287 104
rect 266 100 270 102
rect 266 98 267 100
rect 269 98 270 100
rect 266 93 270 98
rect 256 90 261 92
rect 298 99 302 118
rect 321 114 326 123
rect 338 127 350 131
rect 338 125 346 127
rect 348 125 350 127
rect 321 113 335 114
rect 321 111 329 113
rect 331 111 332 113
rect 334 111 335 113
rect 321 110 335 111
rect 300 97 302 99
rect 298 92 302 97
rect 314 105 327 106
rect 314 103 315 105
rect 317 103 319 105
rect 321 103 327 105
rect 314 102 327 103
rect 314 93 318 102
rect 346 109 350 125
rect 346 107 347 109
rect 349 107 350 109
rect 346 105 350 107
rect 345 103 350 105
rect 345 101 346 103
rect 348 101 350 103
rect 345 96 350 101
rect 300 90 302 92
rect 289 89 302 90
rect 289 87 290 89
rect 292 87 302 89
rect 289 86 302 87
rect 298 85 302 86
rect 345 94 346 96
rect 348 94 350 96
rect 345 92 350 94
rect 364 129 369 131
rect 364 127 366 129
rect 368 127 369 129
rect 364 125 369 127
rect 364 121 368 125
rect 364 119 365 121
rect 367 119 368 121
rect 364 103 368 119
rect 443 129 449 130
rect 443 127 444 129
rect 446 127 449 129
rect 443 126 449 127
rect 364 101 369 103
rect 364 99 366 101
rect 368 99 369 101
rect 364 94 369 99
rect 392 113 400 115
rect 412 114 416 123
rect 392 111 393 113
rect 395 111 400 113
rect 392 109 400 111
rect 410 113 425 114
rect 410 111 412 113
rect 414 111 415 113
rect 417 111 419 113
rect 421 111 425 113
rect 410 110 425 111
rect 395 106 400 109
rect 445 113 449 126
rect 445 111 446 113
rect 448 111 449 113
rect 395 105 433 106
rect 395 103 408 105
rect 410 103 433 105
rect 395 102 433 103
rect 445 106 449 111
rect 443 104 449 106
rect 443 102 444 104
rect 446 102 449 104
rect 443 97 449 102
rect 443 95 444 97
rect 446 95 449 97
rect 364 92 366 94
rect 368 92 369 94
rect 364 90 369 92
rect 443 93 449 95
rect 453 129 459 130
rect 453 127 456 129
rect 458 127 459 129
rect 453 126 459 127
rect 533 129 540 131
rect 533 127 534 129
rect 536 127 540 129
rect 453 106 457 126
rect 486 121 490 123
rect 486 119 487 121
rect 489 119 490 121
rect 453 104 459 106
rect 453 102 456 104
rect 458 102 459 104
rect 453 100 459 102
rect 453 98 456 100
rect 458 98 459 100
rect 453 97 459 98
rect 453 95 456 97
rect 458 95 459 97
rect 453 93 459 95
rect 486 114 490 119
rect 533 125 537 127
rect 539 125 540 127
rect 534 124 540 125
rect 477 113 492 114
rect 477 111 481 113
rect 483 111 488 113
rect 490 111 492 113
rect 477 110 492 111
rect 502 113 510 115
rect 502 111 507 113
rect 509 111 510 113
rect 502 109 510 111
rect 502 108 507 109
rect 502 106 504 108
rect 506 106 507 108
rect 469 102 507 106
rect 534 103 538 124
rect 543 119 547 120
rect 543 117 544 119
rect 546 117 547 119
rect 543 114 547 117
rect 543 113 564 114
rect 543 111 558 113
rect 560 111 564 113
rect 543 110 564 111
rect 574 122 579 124
rect 574 120 575 122
rect 577 120 579 122
rect 574 118 579 120
rect 533 101 538 103
rect 533 99 534 101
rect 536 99 538 101
rect 533 94 538 99
rect 533 92 534 94
rect 536 92 538 94
rect 543 104 548 106
rect 550 104 564 106
rect 543 102 564 104
rect 543 100 547 102
rect 543 98 544 100
rect 546 98 547 100
rect 543 93 547 98
rect 533 90 538 92
rect 575 99 579 118
rect 598 114 603 123
rect 615 127 627 131
rect 615 125 623 127
rect 625 125 627 127
rect 598 113 612 114
rect 598 111 606 113
rect 608 111 609 113
rect 611 111 612 113
rect 598 110 612 111
rect 577 97 579 99
rect 575 92 579 97
rect 591 105 604 106
rect 591 103 592 105
rect 594 103 596 105
rect 598 103 604 105
rect 591 102 604 103
rect 591 93 595 102
rect 623 109 627 125
rect 623 107 624 109
rect 626 107 627 109
rect 623 105 627 107
rect 622 103 627 105
rect 622 101 623 103
rect 625 101 627 103
rect 622 96 627 101
rect 577 90 579 92
rect 566 89 579 90
rect 566 87 567 89
rect 569 87 579 89
rect 566 86 579 87
rect 575 85 579 86
rect 622 94 623 96
rect 625 94 627 96
rect 622 92 627 94
rect 640 129 645 131
rect 640 127 642 129
rect 644 127 645 129
rect 640 125 645 127
rect 640 121 644 125
rect 640 119 641 121
rect 643 119 644 121
rect 640 103 644 119
rect 719 129 725 130
rect 719 127 720 129
rect 722 127 725 129
rect 719 126 725 127
rect 640 101 645 103
rect 640 99 642 101
rect 644 99 645 101
rect 640 94 645 99
rect 668 113 676 115
rect 688 114 692 123
rect 668 111 669 113
rect 671 111 676 113
rect 668 109 676 111
rect 686 113 701 114
rect 686 111 688 113
rect 690 111 691 113
rect 693 111 695 113
rect 697 111 701 113
rect 686 110 701 111
rect 671 106 676 109
rect 721 113 725 126
rect 721 111 722 113
rect 724 111 725 113
rect 671 105 709 106
rect 671 103 684 105
rect 686 103 709 105
rect 671 102 709 103
rect 721 106 725 111
rect 719 104 725 106
rect 719 102 720 104
rect 722 102 725 104
rect 719 97 725 102
rect 719 95 720 97
rect 722 95 725 97
rect 640 92 642 94
rect 644 92 645 94
rect 640 90 645 92
rect 719 93 725 95
rect 729 129 735 130
rect 729 127 732 129
rect 734 127 735 129
rect 729 126 735 127
rect 809 129 816 131
rect 809 127 810 129
rect 812 127 816 129
rect 729 106 733 126
rect 762 121 766 123
rect 762 119 763 121
rect 765 119 766 121
rect 729 104 735 106
rect 729 102 732 104
rect 734 102 735 104
rect 729 100 735 102
rect 729 98 732 100
rect 734 98 735 100
rect 729 97 735 98
rect 729 95 732 97
rect 734 95 735 97
rect 729 93 735 95
rect 762 114 766 119
rect 809 125 813 127
rect 815 125 816 127
rect 810 124 816 125
rect 753 113 768 114
rect 753 111 757 113
rect 759 111 764 113
rect 766 111 768 113
rect 753 110 768 111
rect 778 113 786 115
rect 778 111 783 113
rect 785 111 786 113
rect 778 109 786 111
rect 778 108 783 109
rect 778 106 780 108
rect 782 106 783 108
rect 745 102 783 106
rect 810 103 814 124
rect 819 119 823 120
rect 819 117 820 119
rect 822 117 823 119
rect 819 114 823 117
rect 819 113 840 114
rect 819 111 834 113
rect 836 111 840 113
rect 819 110 840 111
rect 850 122 855 124
rect 850 120 851 122
rect 853 120 855 122
rect 850 118 855 120
rect 809 101 814 103
rect 809 99 810 101
rect 812 99 814 101
rect 809 94 814 99
rect 809 92 810 94
rect 812 92 814 94
rect 819 104 824 106
rect 826 104 840 106
rect 819 102 840 104
rect 819 100 823 102
rect 819 98 820 100
rect 822 98 823 100
rect 819 93 823 98
rect 809 90 814 92
rect 851 99 855 118
rect 874 114 879 123
rect 891 127 903 131
rect 891 125 899 127
rect 901 125 903 127
rect 874 113 888 114
rect 874 111 882 113
rect 884 111 885 113
rect 887 111 888 113
rect 874 110 888 111
rect 853 97 855 99
rect 851 92 855 97
rect 867 105 880 106
rect 867 103 868 105
rect 870 103 872 105
rect 874 103 880 105
rect 867 102 880 103
rect 867 93 871 102
rect 899 109 903 125
rect 899 107 900 109
rect 902 107 903 109
rect 899 105 903 107
rect 898 103 903 105
rect 898 101 899 103
rect 901 101 903 103
rect 898 96 903 101
rect 853 90 855 92
rect 842 89 855 90
rect 842 87 843 89
rect 845 87 855 89
rect 842 86 855 87
rect 851 85 855 86
rect 898 94 899 96
rect 901 94 903 96
rect 898 92 903 94
rect 917 129 922 131
rect 917 127 919 129
rect 921 127 922 129
rect 917 125 922 127
rect 917 121 921 125
rect 917 119 918 121
rect 920 119 921 121
rect 917 103 921 119
rect 996 129 1002 130
rect 996 127 997 129
rect 999 127 1002 129
rect 996 126 1002 127
rect 917 101 922 103
rect 917 99 919 101
rect 921 99 922 101
rect 917 94 922 99
rect 945 113 953 115
rect 965 114 969 123
rect 945 111 946 113
rect 948 111 953 113
rect 945 109 953 111
rect 963 113 978 114
rect 963 111 965 113
rect 967 111 968 113
rect 970 111 972 113
rect 974 111 978 113
rect 963 110 978 111
rect 948 106 953 109
rect 998 113 1002 126
rect 998 111 999 113
rect 1001 111 1002 113
rect 948 105 986 106
rect 948 103 961 105
rect 963 103 986 105
rect 948 102 986 103
rect 998 106 1002 111
rect 996 104 1002 106
rect 996 102 997 104
rect 999 102 1002 104
rect 996 97 1002 102
rect 996 95 997 97
rect 999 95 1002 97
rect 917 92 919 94
rect 921 92 922 94
rect 917 90 922 92
rect 996 93 1002 95
rect 1006 129 1012 130
rect 1006 127 1009 129
rect 1011 127 1012 129
rect 1006 126 1012 127
rect 1086 129 1093 131
rect 1086 127 1087 129
rect 1089 127 1090 129
rect 1092 127 1093 129
rect 1006 106 1010 126
rect 1039 121 1043 123
rect 1039 119 1040 121
rect 1042 119 1043 121
rect 1006 104 1012 106
rect 1006 102 1009 104
rect 1011 102 1012 104
rect 1006 100 1012 102
rect 1006 98 1009 100
rect 1011 98 1012 100
rect 1006 97 1012 98
rect 1006 95 1009 97
rect 1011 95 1012 97
rect 1006 93 1012 95
rect 1039 114 1043 119
rect 1086 125 1093 127
rect 1087 124 1093 125
rect 1030 113 1045 114
rect 1030 111 1034 113
rect 1036 111 1041 113
rect 1043 111 1045 113
rect 1030 110 1045 111
rect 1055 113 1063 115
rect 1055 111 1060 113
rect 1062 111 1063 113
rect 1055 109 1063 111
rect 1055 108 1060 109
rect 1055 106 1057 108
rect 1059 106 1060 108
rect 1022 102 1060 106
rect 1087 103 1091 124
rect 1096 119 1100 120
rect 1096 117 1097 119
rect 1099 117 1100 119
rect 1096 114 1100 117
rect 1096 113 1117 114
rect 1096 111 1111 113
rect 1113 111 1117 113
rect 1096 110 1117 111
rect 1127 122 1132 124
rect 1127 120 1128 122
rect 1130 120 1132 122
rect 1127 118 1132 120
rect 1086 101 1091 103
rect 1086 99 1087 101
rect 1089 99 1091 101
rect 1086 94 1091 99
rect 1086 92 1087 94
rect 1089 92 1091 94
rect 1096 104 1101 106
rect 1103 104 1117 106
rect 1096 102 1117 104
rect 1096 100 1100 102
rect 1096 98 1097 100
rect 1099 98 1100 100
rect 1096 93 1100 98
rect 1086 90 1091 92
rect 1128 99 1132 118
rect 1130 97 1132 99
rect 1128 92 1132 97
rect 1130 90 1132 92
rect 1119 89 1132 90
rect 1119 87 1120 89
rect 1122 87 1132 89
rect 1119 86 1132 87
rect 1128 85 1132 86
rect -287 79 1136 80
rect -287 77 -247 79
rect -245 77 -5 79
rect -3 77 38 79
rect 40 77 78 79
rect 80 77 297 79
rect 299 77 345 79
rect 347 77 574 79
rect 576 77 622 79
rect 624 77 850 79
rect 852 77 898 79
rect 900 77 1127 79
rect 1129 77 1136 79
rect -287 74 1136 77
rect -287 73 1069 74
rect -287 71 99 73
rect 101 72 1069 73
rect 1071 72 1136 74
rect 101 71 1136 72
rect -287 67 1136 71
rect -287 65 -247 67
rect -245 65 -5 67
rect -3 65 38 67
rect 40 65 78 67
rect 80 65 297 67
rect 299 65 345 67
rect 347 65 574 67
rect 576 65 622 67
rect 624 65 850 67
rect 852 65 898 67
rect 900 65 1127 67
rect 1129 65 1136 67
rect -287 64 1136 65
rect -283 58 -271 59
rect -290 54 -271 58
rect -283 53 -271 54
rect -283 51 -282 53
rect -280 51 -278 53
rect -283 41 -278 51
rect -4 58 0 59
rect -13 54 0 58
rect -215 52 -210 54
rect -283 39 -281 41
rect -279 39 -278 41
rect -283 37 -278 39
rect -267 33 -262 35
rect -267 31 -265 33
rect -263 31 -262 33
rect -267 28 -262 31
rect -239 50 -223 51
rect -239 48 -237 50
rect -235 48 -223 50
rect -239 46 -223 48
rect -227 34 -223 46
rect -227 32 -226 34
rect -224 32 -223 34
rect -267 27 -265 28
rect -275 26 -265 27
rect -263 26 -262 28
rect -275 21 -262 26
rect -227 18 -223 32
rect -247 17 -223 18
rect -247 15 -245 17
rect -243 15 -223 17
rect -247 14 -223 15
rect -215 50 -213 52
rect -211 50 -210 52
rect -215 45 -210 50
rect -215 43 -213 45
rect -211 43 -210 45
rect -215 41 -210 43
rect -215 25 -211 41
rect -184 38 -146 42
rect -184 35 -179 38
rect -187 34 -179 35
rect -187 33 -182 34
rect -187 31 -186 33
rect -184 32 -182 33
rect -180 32 -179 34
rect -184 31 -179 32
rect -187 29 -179 31
rect -169 33 -154 34
rect -169 31 -167 33
rect -165 31 -163 33
rect -161 31 -160 33
rect -158 31 -154 33
rect -169 30 -154 31
rect -215 23 -214 25
rect -212 23 -211 25
rect -215 19 -211 23
rect -215 17 -210 19
rect -167 21 -163 30
rect -136 49 -130 51
rect -136 47 -135 49
rect -133 47 -130 49
rect -136 42 -130 47
rect -136 40 -135 42
rect -133 40 -130 42
rect -136 38 -130 40
rect -134 33 -130 38
rect -134 31 -133 33
rect -131 31 -130 33
rect -134 18 -130 31
rect -215 15 -213 17
rect -211 15 -210 17
rect -215 13 -210 15
rect -136 17 -130 18
rect -136 15 -135 17
rect -133 15 -130 17
rect -136 14 -130 15
rect -126 49 -120 51
rect -46 52 -41 54
rect -46 50 -45 52
rect -43 50 -41 52
rect -126 47 -123 49
rect -121 47 -120 49
rect -126 46 -120 47
rect -126 44 -123 46
rect -121 44 -120 46
rect -126 42 -120 44
rect -126 40 -123 42
rect -121 40 -120 42
rect -126 38 -120 40
rect -126 18 -122 38
rect -110 41 -72 42
rect -110 39 -88 41
rect -86 39 -72 41
rect -110 38 -72 39
rect -77 35 -72 38
rect -102 33 -87 34
rect -102 31 -98 33
rect -96 31 -91 33
rect -89 31 -87 33
rect -102 30 -87 31
rect -77 33 -69 35
rect -77 31 -72 33
rect -70 31 -69 33
rect -93 25 -89 30
rect -77 29 -69 31
rect -46 45 -41 50
rect -46 43 -45 45
rect -43 43 -41 45
rect -46 41 -41 43
rect -93 23 -92 25
rect -90 23 -89 25
rect -93 21 -89 23
rect -126 17 -120 18
rect -126 15 -123 17
rect -121 15 -120 17
rect -126 14 -120 15
rect -45 22 -41 41
rect -36 46 -32 51
rect -36 44 -35 46
rect -33 44 -32 46
rect -36 42 -32 44
rect -36 40 -15 42
rect -36 38 -31 40
rect -29 38 -15 40
rect -45 20 -44 22
rect -42 20 -41 22
rect -36 33 -15 34
rect -36 31 -35 33
rect -33 31 -21 33
rect -19 31 -15 33
rect -36 30 -15 31
rect -2 52 0 54
rect -4 47 0 52
rect -2 45 0 47
rect -36 21 -32 30
rect -4 31 0 45
rect 7 44 11 51
rect 38 50 43 52
rect 7 42 8 44
rect 10 42 11 44
rect 7 41 20 42
rect 7 39 12 41
rect 14 39 20 41
rect 7 38 20 39
rect -4 29 -3 31
rect -1 29 0 31
rect -4 26 0 29
rect -5 24 0 26
rect -5 22 -4 24
rect -2 22 0 24
rect -5 20 0 22
rect 14 33 28 34
rect 14 31 22 33
rect 24 31 28 33
rect 14 30 28 31
rect 38 48 39 50
rect 41 48 43 50
rect 38 43 43 48
rect 38 41 39 43
rect 41 41 43 43
rect 38 39 43 41
rect 14 24 19 30
rect 14 22 15 24
rect 17 22 19 24
rect 14 21 19 22
rect -45 19 -41 20
rect -46 17 -41 19
rect 39 19 43 39
rect 47 50 51 51
rect 47 48 48 50
rect 50 48 51 50
rect 47 42 51 48
rect 298 58 302 59
rect 289 54 302 58
rect 87 52 92 54
rect 78 50 83 52
rect 47 41 60 42
rect 47 39 52 41
rect 54 39 60 41
rect 47 38 60 39
rect 54 33 68 34
rect 54 31 62 33
rect 64 31 68 33
rect 54 30 68 31
rect 78 48 79 50
rect 81 48 83 50
rect 78 43 83 48
rect 78 41 79 43
rect 81 41 83 43
rect 78 39 83 41
rect 54 27 59 30
rect 54 25 56 27
rect 58 25 59 27
rect 54 21 59 25
rect 79 33 83 39
rect 79 31 80 33
rect 82 31 83 33
rect -46 15 -45 17
rect -43 15 -41 17
rect -46 13 -41 15
rect 31 17 39 19
rect 41 17 43 19
rect 79 19 83 31
rect 31 15 32 17
rect 34 15 43 17
rect 31 13 43 15
rect 71 17 79 19
rect 81 17 83 19
rect 71 13 83 17
rect 87 50 89 52
rect 91 50 92 52
rect 87 45 92 50
rect 87 43 89 45
rect 91 43 92 45
rect 87 41 92 43
rect 87 25 91 41
rect 118 41 156 42
rect 118 39 133 41
rect 135 39 156 41
rect 118 38 156 39
rect 118 35 123 38
rect 115 33 123 35
rect 115 31 116 33
rect 118 31 123 33
rect 115 29 123 31
rect 133 33 148 34
rect 133 31 135 33
rect 137 31 138 33
rect 140 31 142 33
rect 144 31 148 33
rect 133 30 148 31
rect 87 23 88 25
rect 90 23 91 25
rect 87 19 91 23
rect 87 17 92 19
rect 135 21 139 30
rect 166 49 172 51
rect 166 47 167 49
rect 169 47 172 49
rect 166 42 172 47
rect 166 40 167 42
rect 169 40 172 42
rect 166 38 172 40
rect 168 33 172 38
rect 168 31 169 33
rect 171 31 172 33
rect 168 18 172 31
rect 87 15 89 17
rect 91 15 92 17
rect 87 13 92 15
rect 166 17 172 18
rect 166 15 167 17
rect 169 15 172 17
rect 166 14 172 15
rect 176 49 182 51
rect 256 52 261 54
rect 256 50 257 52
rect 259 50 261 52
rect 176 47 179 49
rect 181 47 182 49
rect 176 46 182 47
rect 176 44 179 46
rect 181 44 182 46
rect 176 42 182 44
rect 176 40 179 42
rect 181 40 182 42
rect 176 38 182 40
rect 176 18 180 38
rect 192 41 230 42
rect 192 39 226 41
rect 228 39 230 41
rect 192 38 230 39
rect 225 35 230 38
rect 200 33 215 34
rect 200 31 204 33
rect 206 31 211 33
rect 213 31 215 33
rect 200 30 215 31
rect 225 33 233 35
rect 225 31 230 33
rect 232 31 233 33
rect 209 25 213 30
rect 225 29 233 31
rect 256 45 261 50
rect 256 43 257 45
rect 259 43 261 45
rect 256 41 261 43
rect 209 23 210 25
rect 212 23 213 25
rect 209 21 213 23
rect 176 17 182 18
rect 176 15 179 17
rect 181 15 182 17
rect 176 14 182 15
rect 257 23 261 41
rect 266 50 270 51
rect 266 48 267 50
rect 269 48 270 50
rect 266 42 270 48
rect 266 40 287 42
rect 266 38 271 40
rect 273 38 287 40
rect 257 21 258 23
rect 260 21 261 23
rect 266 33 287 34
rect 266 31 267 33
rect 269 31 281 33
rect 283 31 287 33
rect 266 30 287 31
rect 300 52 302 54
rect 298 47 302 52
rect 300 45 302 47
rect 266 21 270 30
rect 298 33 302 45
rect 314 49 318 51
rect 314 47 315 49
rect 317 47 318 49
rect 314 42 318 47
rect 575 58 579 59
rect 566 54 579 58
rect 364 52 369 54
rect 345 50 350 52
rect 314 41 327 42
rect 314 39 319 41
rect 321 39 327 41
rect 314 38 327 39
rect 298 31 299 33
rect 301 31 302 33
rect 298 26 302 31
rect 297 24 302 26
rect 297 22 298 24
rect 300 22 302 24
rect 257 19 261 21
rect 297 20 302 22
rect 321 33 335 34
rect 321 31 329 33
rect 331 31 332 33
rect 334 31 335 33
rect 321 30 335 31
rect 345 48 346 50
rect 348 48 350 50
rect 345 43 350 48
rect 345 41 346 43
rect 348 41 350 43
rect 345 39 350 41
rect 321 21 326 30
rect 346 37 347 39
rect 349 37 350 39
rect 256 17 261 19
rect 346 19 350 37
rect 256 15 257 17
rect 259 15 261 17
rect 256 13 261 15
rect 338 17 346 19
rect 348 17 350 19
rect 338 13 350 17
rect 364 50 366 52
rect 368 50 369 52
rect 364 45 369 50
rect 364 43 366 45
rect 368 43 369 45
rect 364 41 369 43
rect 364 25 368 41
rect 395 41 433 42
rect 395 39 410 41
rect 412 39 433 41
rect 395 38 433 39
rect 395 35 400 38
rect 392 33 400 35
rect 392 31 393 33
rect 395 31 400 33
rect 392 29 400 31
rect 410 33 425 34
rect 410 31 412 33
rect 414 31 415 33
rect 417 31 419 33
rect 421 31 425 33
rect 410 30 425 31
rect 364 23 365 25
rect 367 23 368 25
rect 364 19 368 23
rect 364 17 369 19
rect 412 21 416 30
rect 443 49 449 51
rect 443 47 444 49
rect 446 47 449 49
rect 443 42 449 47
rect 443 40 444 42
rect 446 40 449 42
rect 443 38 449 40
rect 445 33 449 38
rect 445 31 446 33
rect 448 31 449 33
rect 445 18 449 31
rect 364 15 366 17
rect 368 15 369 17
rect 364 13 369 15
rect 443 17 449 18
rect 443 15 444 17
rect 446 15 449 17
rect 443 14 449 15
rect 453 49 459 51
rect 533 52 538 54
rect 533 50 534 52
rect 536 50 538 52
rect 453 47 456 49
rect 458 47 459 49
rect 453 46 459 47
rect 453 44 456 46
rect 458 44 459 46
rect 453 42 459 44
rect 453 40 456 42
rect 458 40 459 42
rect 453 38 459 40
rect 453 18 457 38
rect 469 41 507 42
rect 469 39 503 41
rect 505 39 507 41
rect 469 38 507 39
rect 502 35 507 38
rect 477 33 492 34
rect 477 31 481 33
rect 483 31 488 33
rect 490 31 492 33
rect 477 30 492 31
rect 502 33 510 35
rect 502 31 507 33
rect 509 31 510 33
rect 486 25 490 30
rect 502 29 510 31
rect 533 45 538 50
rect 533 43 534 45
rect 536 43 538 45
rect 533 41 538 43
rect 486 23 487 25
rect 489 23 490 25
rect 486 21 490 23
rect 453 17 459 18
rect 453 15 456 17
rect 458 15 459 17
rect 453 14 459 15
rect 534 23 538 41
rect 543 50 547 51
rect 543 48 544 50
rect 546 48 547 50
rect 543 42 547 48
rect 543 40 564 42
rect 543 38 548 40
rect 550 38 564 40
rect 534 21 535 23
rect 537 21 538 23
rect 543 33 564 34
rect 543 31 544 33
rect 546 31 558 33
rect 560 31 564 33
rect 543 30 564 31
rect 577 52 579 54
rect 575 47 579 52
rect 577 45 579 47
rect 543 21 547 30
rect 575 33 579 45
rect 591 49 595 51
rect 591 47 592 49
rect 594 47 595 49
rect 591 42 595 47
rect 851 58 855 59
rect 842 54 855 58
rect 640 52 645 54
rect 622 50 627 52
rect 591 41 604 42
rect 591 39 596 41
rect 598 39 604 41
rect 591 38 604 39
rect 575 31 576 33
rect 578 31 579 33
rect 575 26 579 31
rect 574 24 579 26
rect 574 22 575 24
rect 577 22 579 24
rect 534 19 538 21
rect 574 20 579 22
rect 598 33 612 34
rect 598 31 606 33
rect 608 31 609 33
rect 611 31 612 33
rect 598 30 612 31
rect 622 48 623 50
rect 625 48 627 50
rect 622 43 627 48
rect 622 41 623 43
rect 625 41 627 43
rect 622 39 627 41
rect 598 21 603 30
rect 623 37 624 39
rect 626 37 627 39
rect 533 17 538 19
rect 623 19 627 37
rect 533 15 534 17
rect 536 15 538 17
rect 533 13 538 15
rect 615 17 623 19
rect 625 17 627 19
rect 615 13 627 17
rect 640 50 642 52
rect 644 50 645 52
rect 640 45 645 50
rect 640 43 642 45
rect 644 43 645 45
rect 640 41 645 43
rect 640 25 644 41
rect 671 41 709 42
rect 671 39 686 41
rect 688 39 709 41
rect 671 38 709 39
rect 671 35 676 38
rect 668 33 676 35
rect 668 31 669 33
rect 671 31 676 33
rect 668 29 676 31
rect 686 33 701 34
rect 686 31 688 33
rect 690 31 691 33
rect 693 31 695 33
rect 697 31 701 33
rect 686 30 701 31
rect 640 23 641 25
rect 643 23 644 25
rect 640 19 644 23
rect 640 17 645 19
rect 688 21 692 30
rect 719 49 725 51
rect 719 47 720 49
rect 722 47 725 49
rect 719 42 725 47
rect 719 40 720 42
rect 722 40 725 42
rect 719 38 725 40
rect 721 33 725 38
rect 721 31 722 33
rect 724 31 725 33
rect 721 18 725 31
rect 640 15 642 17
rect 644 15 645 17
rect 640 13 645 15
rect 719 17 725 18
rect 719 15 720 17
rect 722 15 725 17
rect 719 14 725 15
rect 729 49 735 51
rect 809 52 814 54
rect 809 50 810 52
rect 812 50 814 52
rect 729 47 732 49
rect 734 47 735 49
rect 729 46 735 47
rect 729 44 732 46
rect 734 44 735 46
rect 729 42 735 44
rect 729 40 732 42
rect 734 40 735 42
rect 729 38 735 40
rect 729 18 733 38
rect 745 41 783 42
rect 745 39 779 41
rect 781 39 783 41
rect 745 38 783 39
rect 778 35 783 38
rect 753 33 768 34
rect 753 31 757 33
rect 759 31 764 33
rect 766 31 768 33
rect 753 30 768 31
rect 778 33 786 35
rect 778 31 783 33
rect 785 31 786 33
rect 762 25 766 30
rect 778 29 786 31
rect 809 45 814 50
rect 809 43 810 45
rect 812 43 814 45
rect 809 41 814 43
rect 762 23 763 25
rect 765 23 766 25
rect 762 21 766 23
rect 729 17 735 18
rect 729 15 732 17
rect 734 15 735 17
rect 729 14 735 15
rect 810 23 814 41
rect 819 50 823 51
rect 819 48 820 50
rect 822 48 823 50
rect 819 42 823 48
rect 819 40 840 42
rect 819 38 824 40
rect 826 38 840 40
rect 810 21 811 23
rect 813 21 814 23
rect 819 33 840 34
rect 819 31 820 33
rect 822 31 834 33
rect 836 31 840 33
rect 819 30 840 31
rect 853 52 855 54
rect 851 47 855 52
rect 853 45 855 47
rect 819 21 823 30
rect 851 33 855 45
rect 867 49 871 51
rect 867 47 868 49
rect 870 47 871 49
rect 867 42 871 47
rect 1128 58 1132 59
rect 1119 54 1132 58
rect 917 52 922 54
rect 898 50 903 52
rect 867 41 880 42
rect 867 39 872 41
rect 874 39 880 41
rect 867 38 880 39
rect 851 31 852 33
rect 854 31 855 33
rect 851 26 855 31
rect 850 24 855 26
rect 850 22 851 24
rect 853 22 855 24
rect 810 19 814 21
rect 850 20 855 22
rect 874 33 888 34
rect 874 31 882 33
rect 884 31 885 33
rect 887 31 888 33
rect 874 30 888 31
rect 898 48 899 50
rect 901 48 903 50
rect 898 43 903 48
rect 898 41 899 43
rect 901 41 903 43
rect 898 39 903 41
rect 874 21 879 30
rect 899 37 900 39
rect 902 37 903 39
rect 809 17 814 19
rect 899 19 903 37
rect 809 15 810 17
rect 812 15 814 17
rect 809 13 814 15
rect 891 17 899 19
rect 901 17 903 19
rect 891 13 903 17
rect 917 50 919 52
rect 921 50 922 52
rect 917 45 922 50
rect 917 43 919 45
rect 921 43 922 45
rect 917 41 922 43
rect 917 25 921 41
rect 948 41 986 42
rect 948 39 963 41
rect 965 39 986 41
rect 948 38 986 39
rect 948 35 953 38
rect 945 33 953 35
rect 945 31 946 33
rect 948 31 953 33
rect 945 29 953 31
rect 963 33 978 34
rect 963 31 965 33
rect 967 31 968 33
rect 970 31 972 33
rect 974 31 978 33
rect 963 30 978 31
rect 917 23 918 25
rect 920 23 921 25
rect 917 19 921 23
rect 917 17 922 19
rect 965 21 969 30
rect 996 49 1002 51
rect 996 47 997 49
rect 999 47 1002 49
rect 996 42 1002 47
rect 996 40 997 42
rect 999 40 1002 42
rect 996 38 1002 40
rect 998 33 1002 38
rect 998 31 999 33
rect 1001 31 1002 33
rect 998 18 1002 31
rect 917 15 919 17
rect 921 15 922 17
rect 917 13 922 15
rect 996 17 1002 18
rect 996 15 997 17
rect 999 15 1002 17
rect 996 14 1002 15
rect 1006 49 1012 51
rect 1086 52 1091 54
rect 1086 50 1087 52
rect 1089 50 1091 52
rect 1006 47 1009 49
rect 1011 47 1012 49
rect 1006 46 1012 47
rect 1006 44 1009 46
rect 1011 44 1012 46
rect 1006 42 1012 44
rect 1006 40 1009 42
rect 1011 40 1012 42
rect 1006 38 1012 40
rect 1006 18 1010 38
rect 1022 41 1060 42
rect 1022 39 1056 41
rect 1058 39 1060 41
rect 1022 38 1060 39
rect 1055 35 1060 38
rect 1030 33 1045 34
rect 1030 31 1034 33
rect 1036 31 1041 33
rect 1043 31 1045 33
rect 1030 30 1045 31
rect 1055 33 1063 35
rect 1055 31 1060 33
rect 1062 31 1063 33
rect 1039 25 1043 30
rect 1055 29 1063 31
rect 1086 45 1091 50
rect 1086 43 1087 45
rect 1089 43 1091 45
rect 1086 41 1091 43
rect 1039 23 1040 25
rect 1042 23 1043 25
rect 1039 21 1043 23
rect 1006 17 1012 18
rect 1006 15 1009 17
rect 1011 15 1012 17
rect 1006 14 1012 15
rect 1087 20 1091 41
rect 1096 50 1100 51
rect 1096 48 1097 50
rect 1099 48 1100 50
rect 1096 42 1100 48
rect 1096 40 1117 42
rect 1096 38 1101 40
rect 1103 38 1117 40
rect 1096 33 1117 34
rect 1096 31 1097 33
rect 1099 31 1111 33
rect 1113 31 1117 33
rect 1096 30 1117 31
rect 1130 52 1132 54
rect 1128 47 1132 52
rect 1130 45 1132 47
rect 1096 21 1100 30
rect 1128 30 1132 45
rect 1128 28 1129 30
rect 1131 28 1132 30
rect 1128 26 1132 28
rect 1127 24 1132 26
rect 1127 22 1128 24
rect 1130 22 1132 24
rect 1127 20 1132 22
rect 1087 19 1088 20
rect 1086 18 1088 19
rect 1090 18 1091 20
rect 1086 17 1091 18
rect 1086 15 1087 17
rect 1089 15 1091 17
rect 1086 13 1091 15
rect -287 7 1136 8
rect -287 5 -280 7
rect -278 5 -227 7
rect -225 5 -5 7
rect -3 5 28 7
rect 30 5 38 7
rect 40 5 68 7
rect 70 5 78 7
rect 80 5 297 7
rect 299 5 335 7
rect 337 5 345 7
rect 347 5 574 7
rect 576 5 612 7
rect 614 5 622 7
rect 624 5 850 7
rect 852 5 888 7
rect 890 5 898 7
rect 900 5 1127 7
rect 1129 5 1136 7
rect -287 4 164 5
rect -287 2 134 4
rect 136 3 164 4
rect 166 3 1136 5
rect 136 2 1136 3
rect -287 0 1136 2
rect -158 -4 1133 0
rect -158 -6 -153 -4
rect -151 -6 -142 -4
rect -140 -6 -121 -4
rect -119 -6 -113 -4
rect -111 -6 -101 -4
rect -99 -6 -90 -4
rect -88 -6 -69 -4
rect -67 -6 -61 -4
rect -59 -6 -49 -4
rect -47 -6 -38 -4
rect -36 -6 -17 -4
rect -15 -6 -9 -4
rect -7 -6 3 -4
rect 5 -6 14 -4
rect 16 -6 35 -4
rect 37 -6 43 -4
rect 45 -6 55 -4
rect 57 -6 66 -4
rect 68 -6 87 -4
rect 89 -6 95 -4
rect 97 -6 108 -4
rect 110 -6 119 -4
rect 121 -6 140 -4
rect 142 -6 148 -4
rect 150 -6 165 -4
rect 167 -6 173 -4
rect 175 -6 185 -4
rect 187 -6 193 -4
rect 195 -6 205 -4
rect 207 -6 213 -4
rect 215 -6 227 -4
rect 229 -6 235 -4
rect 237 -6 249 -4
rect 251 -6 257 -4
rect 259 -6 271 -4
rect 273 -6 279 -4
rect 281 -6 296 -4
rect 298 -6 307 -4
rect 309 -6 328 -4
rect 330 -6 336 -4
rect 338 -6 349 -4
rect 351 -6 360 -4
rect 362 -6 381 -4
rect 383 -6 389 -4
rect 391 -6 401 -4
rect 403 -6 412 -4
rect 414 -6 433 -4
rect 435 -6 441 -4
rect 443 -6 453 -4
rect 455 -6 464 -4
rect 466 -6 485 -4
rect 487 -6 493 -4
rect 495 -6 505 -4
rect 507 -6 516 -4
rect 518 -6 537 -4
rect 539 -6 545 -4
rect 547 -6 560 -4
rect 562 -6 568 -4
rect 570 -6 581 -4
rect 583 -6 589 -4
rect 591 -6 604 -4
rect 606 -6 615 -4
rect 617 -6 636 -4
rect 638 -6 644 -4
rect 646 -6 657 -4
rect 659 -6 668 -4
rect 670 -6 689 -4
rect 691 -6 697 -4
rect 699 -6 709 -4
rect 711 -6 720 -4
rect 722 -6 741 -4
rect 743 -6 749 -4
rect 751 -6 761 -4
rect 763 -6 772 -4
rect 774 -6 793 -4
rect 795 -6 801 -4
rect 803 -6 813 -4
rect 815 -6 824 -4
rect 826 -6 845 -4
rect 847 -6 853 -4
rect 855 -6 865 -4
rect 867 -6 876 -4
rect 878 -6 897 -4
rect 899 -6 905 -4
rect 907 -6 918 -4
rect 920 -6 929 -4
rect 931 -6 950 -4
rect 952 -6 958 -4
rect 960 -6 972 -4
rect 974 -6 983 -4
rect 985 -6 1004 -4
rect 1006 -6 1012 -4
rect 1014 -6 1027 -4
rect 1029 -6 1038 -4
rect 1040 -6 1059 -4
rect 1061 -6 1067 -4
rect 1069 -6 1080 -4
rect 1082 -6 1091 -4
rect 1093 -6 1112 -4
rect 1114 -6 1120 -4
rect 1122 -6 1133 -4
rect -158 -7 1133 -6
rect -156 -21 -152 -12
rect -156 -23 -154 -21
rect -156 -52 -152 -23
rect -132 -21 -128 -20
rect -132 -23 -131 -21
rect -129 -23 -128 -21
rect -132 -29 -128 -23
rect -141 -30 -128 -29
rect -141 -32 -137 -30
rect -135 -32 -128 -30
rect -141 -33 -128 -32
rect -124 -29 -120 -20
rect -104 -21 -100 -12
rect -104 -23 -102 -21
rect -124 -30 -111 -29
rect -124 -32 -115 -30
rect -113 -32 -111 -30
rect -124 -33 -111 -32
rect -133 -38 -121 -37
rect -133 -40 -125 -38
rect -123 -40 -121 -38
rect -133 -41 -121 -40
rect -117 -38 -111 -33
rect -117 -40 -114 -38
rect -112 -40 -111 -38
rect -117 -41 -111 -40
rect -125 -45 -121 -41
rect -125 -46 -111 -45
rect -125 -48 -120 -46
rect -118 -48 -111 -46
rect -125 -49 -111 -48
rect -104 -52 -100 -23
rect -80 -21 -76 -20
rect -80 -23 -79 -21
rect -77 -23 -76 -21
rect -80 -29 -76 -23
rect -89 -30 -76 -29
rect -89 -32 -85 -30
rect -83 -32 -76 -30
rect -89 -33 -76 -32
rect -72 -29 -68 -20
rect -52 -21 -48 -12
rect -52 -23 -50 -21
rect -72 -30 -59 -29
rect -72 -32 -63 -30
rect -61 -32 -59 -30
rect -72 -33 -59 -32
rect -81 -38 -69 -37
rect -81 -40 -73 -38
rect -71 -40 -69 -38
rect -81 -41 -69 -40
rect -65 -38 -59 -33
rect -65 -40 -62 -38
rect -60 -40 -59 -38
rect -65 -41 -59 -40
rect -73 -45 -69 -41
rect -73 -46 -59 -45
rect -73 -48 -69 -46
rect -67 -48 -59 -46
rect -73 -49 -59 -48
rect -52 -52 -48 -23
rect -28 -21 -24 -20
rect -28 -23 -27 -21
rect -25 -23 -24 -21
rect -28 -29 -24 -23
rect -37 -30 -24 -29
rect -37 -32 -33 -30
rect -31 -32 -24 -30
rect -37 -33 -24 -32
rect -20 -29 -16 -20
rect 0 -21 4 -12
rect 0 -23 2 -21
rect -20 -30 -7 -29
rect -20 -32 -11 -30
rect -9 -32 -7 -30
rect -20 -33 -7 -32
rect -29 -38 -17 -37
rect -29 -40 -21 -38
rect -19 -40 -17 -38
rect -29 -41 -17 -40
rect -13 -38 -7 -33
rect -13 -40 -10 -38
rect -8 -40 -7 -38
rect -13 -41 -7 -40
rect -21 -45 -17 -41
rect -21 -46 -7 -45
rect -21 -48 -16 -46
rect -14 -48 -7 -46
rect -21 -49 -7 -48
rect 0 -52 4 -23
rect 24 -29 28 -20
rect 15 -30 25 -29
rect 15 -32 19 -30
rect 21 -31 25 -30
rect 27 -31 28 -29
rect 21 -32 28 -31
rect 15 -33 28 -32
rect 32 -29 36 -20
rect 52 -21 56 -12
rect 52 -23 54 -21
rect 32 -30 45 -29
rect 32 -32 41 -30
rect 43 -32 45 -30
rect 32 -33 45 -32
rect 23 -38 35 -37
rect 23 -40 31 -38
rect 33 -40 35 -38
rect 23 -41 35 -40
rect 39 -38 45 -33
rect 39 -40 42 -38
rect 44 -40 45 -38
rect 39 -41 45 -40
rect 31 -45 35 -41
rect 31 -46 45 -45
rect 31 -48 35 -46
rect 37 -48 45 -46
rect 31 -49 45 -48
rect 52 -52 56 -23
rect 76 -27 80 -20
rect 76 -29 77 -27
rect 79 -29 80 -27
rect 67 -30 80 -29
rect 67 -32 71 -30
rect 73 -32 80 -30
rect 67 -33 80 -32
rect 84 -29 88 -20
rect 105 -21 109 -12
rect 105 -23 107 -21
rect 84 -30 97 -29
rect 84 -32 93 -30
rect 95 -32 97 -30
rect 84 -33 97 -32
rect 75 -38 87 -37
rect 75 -40 83 -38
rect 85 -40 87 -38
rect 75 -41 87 -40
rect 91 -38 97 -33
rect 91 -40 94 -38
rect 96 -40 97 -38
rect 91 -41 97 -40
rect 83 -45 87 -41
rect 83 -46 97 -45
rect 83 -48 87 -46
rect 89 -48 97 -46
rect 83 -49 97 -48
rect 105 -52 109 -23
rect 129 -22 133 -20
rect 129 -24 130 -22
rect 132 -24 133 -22
rect 129 -29 133 -24
rect 120 -30 133 -29
rect 120 -32 124 -30
rect 126 -32 133 -30
rect 120 -33 133 -32
rect 137 -29 141 -20
rect 162 -21 168 -20
rect 162 -23 164 -21
rect 166 -23 168 -21
rect 162 -28 168 -23
rect 182 -21 188 -20
rect 182 -23 184 -21
rect 186 -23 188 -21
rect 182 -24 188 -23
rect 202 -21 208 -20
rect 202 -23 204 -21
rect 206 -23 208 -21
rect 182 -26 184 -24
rect 186 -26 188 -24
rect 182 -28 188 -26
rect 202 -28 208 -23
rect 224 -21 230 -20
rect 224 -23 226 -21
rect 228 -23 230 -21
rect 224 -28 230 -23
rect 246 -21 252 -20
rect 246 -23 248 -21
rect 250 -23 252 -21
rect 246 -28 252 -23
rect 268 -21 274 -20
rect 268 -23 270 -21
rect 272 -23 274 -21
rect 268 -28 274 -23
rect 293 -21 297 -12
rect 293 -23 295 -21
rect 137 -30 150 -29
rect 137 -32 146 -30
rect 148 -32 150 -30
rect 137 -33 150 -32
rect 128 -38 140 -37
rect 128 -40 136 -38
rect 138 -40 140 -38
rect 128 -41 140 -40
rect 144 -38 150 -33
rect 162 -34 174 -28
rect 182 -34 194 -28
rect 202 -31 214 -28
rect 202 -33 210 -31
rect 212 -33 214 -31
rect 202 -34 214 -33
rect 224 -31 236 -28
rect 224 -33 230 -31
rect 232 -33 236 -31
rect 224 -34 236 -33
rect 246 -31 258 -28
rect 246 -33 250 -31
rect 252 -33 258 -31
rect 246 -34 258 -33
rect 268 -34 280 -28
rect 144 -40 147 -38
rect 149 -40 150 -38
rect 144 -41 150 -40
rect 170 -38 174 -34
rect 190 -38 194 -34
rect 210 -38 214 -34
rect 232 -38 236 -34
rect 254 -38 258 -34
rect 276 -38 280 -34
rect 170 -40 171 -38
rect 173 -39 178 -38
rect 173 -40 174 -39
rect 170 -41 174 -40
rect 176 -41 178 -39
rect 136 -45 140 -41
rect 170 -42 178 -41
rect 190 -39 198 -38
rect 190 -41 194 -39
rect 196 -41 198 -39
rect 190 -42 198 -41
rect 210 -39 218 -38
rect 210 -41 214 -39
rect 216 -41 218 -39
rect 210 -42 218 -41
rect 232 -39 240 -38
rect 232 -41 236 -39
rect 238 -41 240 -39
rect 232 -42 240 -41
rect 254 -39 262 -38
rect 254 -41 258 -39
rect 260 -41 262 -39
rect 254 -42 262 -41
rect 276 -39 284 -38
rect 276 -41 277 -39
rect 279 -41 280 -39
rect 282 -41 284 -39
rect 276 -42 284 -41
rect 293 -40 297 -23
rect 317 -22 321 -20
rect 317 -24 318 -22
rect 320 -24 321 -22
rect 293 -42 294 -40
rect 296 -42 297 -40
rect 162 -45 166 -44
rect 136 -46 150 -45
rect 136 -48 140 -46
rect 142 -48 150 -46
rect 136 -49 150 -48
rect 162 -47 163 -45
rect 165 -47 166 -45
rect 162 -52 166 -47
rect 182 -45 186 -44
rect 182 -47 183 -45
rect 185 -47 186 -45
rect 182 -52 186 -47
rect 202 -47 206 -44
rect 202 -49 203 -47
rect 205 -49 206 -47
rect 202 -52 206 -49
rect 224 -46 228 -44
rect 224 -48 225 -46
rect 227 -48 228 -46
rect 224 -52 228 -48
rect 246 -48 250 -44
rect 246 -50 247 -48
rect 249 -50 250 -48
rect 246 -52 250 -50
rect 268 -49 272 -44
rect 268 -51 269 -49
rect 271 -51 272 -49
rect 268 -52 272 -51
rect 293 -52 297 -42
rect 317 -29 321 -24
rect 308 -30 321 -29
rect 308 -32 312 -30
rect 314 -32 321 -30
rect 308 -33 321 -32
rect 325 -29 329 -20
rect 346 -21 350 -12
rect 346 -23 348 -21
rect 325 -30 338 -29
rect 325 -32 334 -30
rect 336 -32 338 -30
rect 325 -33 338 -32
rect 316 -38 328 -37
rect 316 -40 324 -38
rect 326 -40 328 -38
rect 316 -41 328 -40
rect 332 -38 338 -33
rect 332 -40 335 -38
rect 337 -40 338 -38
rect 332 -41 338 -40
rect 324 -45 328 -41
rect 324 -46 338 -45
rect 324 -48 329 -46
rect 331 -48 338 -46
rect 324 -49 338 -48
rect 346 -52 350 -23
rect 370 -29 374 -20
rect 361 -30 374 -29
rect 361 -32 365 -30
rect 367 -32 368 -30
rect 370 -32 374 -30
rect 361 -33 374 -32
rect 378 -29 382 -20
rect 398 -21 402 -12
rect 398 -23 400 -21
rect 378 -30 391 -29
rect 378 -32 387 -30
rect 389 -32 391 -30
rect 378 -33 391 -32
rect 369 -38 381 -37
rect 369 -40 377 -38
rect 379 -40 381 -38
rect 369 -41 381 -40
rect 385 -38 391 -33
rect 385 -40 388 -38
rect 390 -40 391 -38
rect 385 -41 391 -40
rect 377 -45 381 -41
rect 377 -46 391 -45
rect 377 -48 382 -46
rect 384 -48 391 -46
rect 377 -49 391 -48
rect 398 -52 402 -23
rect 422 -27 426 -20
rect 422 -29 423 -27
rect 425 -29 426 -27
rect 413 -30 426 -29
rect 413 -32 417 -30
rect 419 -32 426 -30
rect 413 -33 426 -32
rect 430 -29 434 -20
rect 450 -21 454 -12
rect 450 -23 452 -21
rect 430 -30 443 -29
rect 430 -32 439 -30
rect 441 -32 443 -30
rect 430 -33 443 -32
rect 421 -38 433 -37
rect 421 -40 429 -38
rect 431 -40 433 -38
rect 421 -41 433 -40
rect 437 -38 443 -33
rect 437 -40 440 -38
rect 442 -40 443 -38
rect 437 -41 443 -40
rect 429 -45 433 -41
rect 429 -46 443 -45
rect 429 -48 433 -46
rect 435 -48 443 -46
rect 429 -49 443 -48
rect 450 -52 454 -23
rect 474 -29 478 -20
rect 465 -30 478 -29
rect 465 -32 469 -30
rect 471 -32 473 -30
rect 475 -32 478 -30
rect 465 -33 478 -32
rect 482 -29 486 -20
rect 502 -21 506 -12
rect 502 -23 504 -21
rect 482 -30 495 -29
rect 482 -32 491 -30
rect 493 -32 495 -30
rect 482 -33 495 -32
rect 473 -38 485 -37
rect 473 -40 481 -38
rect 483 -40 485 -38
rect 473 -41 485 -40
rect 489 -38 495 -33
rect 489 -40 492 -38
rect 494 -40 495 -38
rect 489 -41 495 -40
rect 481 -45 485 -41
rect 481 -46 495 -45
rect 481 -48 486 -46
rect 488 -48 495 -46
rect 481 -49 495 -48
rect 502 -52 506 -23
rect 526 -26 530 -20
rect 526 -28 527 -26
rect 529 -28 530 -26
rect 526 -29 530 -28
rect 517 -30 530 -29
rect 517 -32 521 -30
rect 523 -32 530 -30
rect 517 -33 530 -32
rect 534 -29 538 -20
rect 557 -21 563 -20
rect 557 -23 559 -21
rect 561 -23 563 -21
rect 557 -28 563 -23
rect 578 -21 584 -20
rect 578 -23 580 -21
rect 582 -23 584 -21
rect 578 -28 584 -23
rect 601 -21 605 -12
rect 601 -23 603 -21
rect 534 -30 547 -29
rect 534 -32 543 -30
rect 545 -32 547 -30
rect 534 -33 547 -32
rect 525 -38 537 -37
rect 525 -40 533 -38
rect 535 -40 537 -38
rect 525 -41 537 -40
rect 541 -38 547 -33
rect 557 -34 569 -28
rect 578 -34 590 -28
rect 541 -40 544 -38
rect 546 -40 547 -38
rect 541 -41 547 -40
rect 565 -36 569 -34
rect 565 -38 566 -36
rect 568 -38 569 -36
rect 586 -38 590 -34
rect 565 -39 573 -38
rect 565 -41 569 -39
rect 571 -41 573 -39
rect 533 -45 537 -41
rect 565 -42 573 -41
rect 586 -40 587 -38
rect 589 -39 594 -38
rect 589 -40 590 -39
rect 586 -41 590 -40
rect 592 -41 594 -39
rect 586 -42 594 -41
rect 533 -46 547 -45
rect 533 -48 537 -46
rect 539 -48 547 -46
rect 533 -49 547 -48
rect 557 -52 561 -44
rect 578 -52 582 -44
rect 601 -52 605 -23
rect 625 -23 629 -20
rect 625 -25 626 -23
rect 628 -25 629 -23
rect 625 -29 629 -25
rect 616 -30 629 -29
rect 616 -32 620 -30
rect 622 -32 629 -30
rect 616 -33 629 -32
rect 633 -29 637 -20
rect 654 -21 658 -12
rect 654 -23 656 -21
rect 633 -30 646 -29
rect 633 -32 642 -30
rect 644 -32 646 -30
rect 633 -33 646 -32
rect 624 -38 636 -37
rect 624 -40 632 -38
rect 634 -40 636 -38
rect 624 -41 636 -40
rect 640 -38 646 -33
rect 640 -40 643 -38
rect 645 -40 646 -38
rect 640 -41 646 -40
rect 632 -45 636 -41
rect 632 -46 646 -45
rect 632 -48 643 -46
rect 645 -48 646 -46
rect 632 -49 646 -48
rect 654 -52 658 -23
rect 678 -21 682 -20
rect 678 -23 679 -21
rect 681 -23 682 -21
rect 678 -29 682 -23
rect 669 -30 682 -29
rect 669 -32 673 -30
rect 675 -32 682 -30
rect 669 -33 682 -32
rect 686 -29 690 -20
rect 706 -21 710 -12
rect 706 -23 708 -21
rect 686 -30 699 -29
rect 686 -32 695 -30
rect 697 -32 699 -30
rect 686 -33 699 -32
rect 677 -38 689 -37
rect 677 -40 685 -38
rect 687 -40 689 -38
rect 677 -41 689 -40
rect 693 -38 699 -33
rect 693 -40 696 -38
rect 698 -40 699 -38
rect 693 -41 699 -40
rect 685 -45 689 -41
rect 685 -46 699 -45
rect 685 -48 690 -46
rect 692 -48 699 -46
rect 685 -49 699 -48
rect 706 -52 710 -23
rect 730 -22 734 -20
rect 730 -24 731 -22
rect 733 -24 734 -22
rect 730 -29 734 -24
rect 721 -30 734 -29
rect 721 -32 725 -30
rect 727 -32 734 -30
rect 721 -33 734 -32
rect 738 -29 742 -20
rect 758 -21 762 -12
rect 758 -23 760 -21
rect 738 -30 751 -29
rect 738 -32 747 -30
rect 749 -32 751 -30
rect 738 -33 751 -32
rect 729 -38 741 -37
rect 729 -40 737 -38
rect 739 -40 741 -38
rect 729 -41 741 -40
rect 745 -38 751 -33
rect 745 -40 748 -38
rect 750 -40 751 -38
rect 745 -41 751 -40
rect 737 -45 741 -41
rect 737 -46 751 -45
rect 737 -48 741 -46
rect 743 -48 751 -46
rect 737 -49 751 -48
rect 758 -52 762 -23
rect 782 -22 786 -20
rect 782 -24 783 -22
rect 785 -24 786 -22
rect 782 -29 786 -24
rect 773 -30 786 -29
rect 773 -32 777 -30
rect 779 -32 786 -30
rect 773 -33 786 -32
rect 790 -29 794 -20
rect 810 -21 814 -12
rect 810 -23 812 -21
rect 790 -30 803 -29
rect 790 -32 799 -30
rect 801 -32 803 -30
rect 790 -33 803 -32
rect 781 -38 793 -37
rect 781 -40 789 -38
rect 791 -40 793 -38
rect 781 -41 793 -40
rect 797 -38 803 -33
rect 797 -40 800 -38
rect 802 -40 803 -38
rect 797 -41 803 -40
rect 789 -45 793 -41
rect 789 -46 803 -45
rect 789 -48 794 -46
rect 796 -48 803 -46
rect 789 -49 803 -48
rect 810 -52 814 -23
rect 834 -22 838 -20
rect 834 -24 835 -22
rect 837 -24 838 -22
rect 834 -29 838 -24
rect 825 -30 838 -29
rect 825 -32 829 -30
rect 831 -32 838 -30
rect 825 -33 838 -32
rect 842 -29 846 -20
rect 862 -21 866 -12
rect 862 -23 864 -21
rect 842 -30 855 -29
rect 842 -32 851 -30
rect 853 -32 855 -30
rect 842 -33 855 -32
rect 833 -38 845 -37
rect 833 -40 841 -38
rect 843 -40 845 -38
rect 833 -41 845 -40
rect 849 -38 855 -33
rect 849 -40 852 -38
rect 854 -40 855 -38
rect 849 -41 855 -40
rect 841 -45 845 -41
rect 841 -46 855 -45
rect 841 -48 845 -46
rect 847 -48 855 -46
rect 841 -49 855 -48
rect 862 -52 866 -23
rect 886 -22 890 -20
rect 886 -24 887 -22
rect 889 -24 890 -22
rect 886 -29 890 -24
rect 877 -30 890 -29
rect 877 -32 881 -30
rect 883 -32 890 -30
rect 877 -33 890 -32
rect 894 -29 898 -20
rect 915 -21 919 -12
rect 915 -23 917 -21
rect 894 -30 907 -29
rect 894 -32 903 -30
rect 905 -32 907 -30
rect 894 -33 907 -32
rect 885 -38 897 -37
rect 885 -40 893 -38
rect 895 -40 897 -38
rect 885 -41 897 -40
rect 901 -38 907 -33
rect 901 -40 904 -38
rect 906 -40 907 -38
rect 901 -41 907 -40
rect 893 -45 897 -41
rect 893 -46 907 -45
rect 893 -48 897 -46
rect 899 -48 907 -46
rect 893 -49 907 -48
rect 915 -52 919 -23
rect 939 -22 943 -20
rect 939 -24 940 -22
rect 942 -24 943 -22
rect 939 -29 943 -24
rect 930 -30 943 -29
rect 930 -32 934 -30
rect 936 -32 943 -30
rect 930 -33 943 -32
rect 947 -29 951 -20
rect 969 -21 973 -12
rect 969 -23 971 -21
rect 947 -30 960 -29
rect 947 -32 956 -30
rect 958 -32 960 -30
rect 947 -33 960 -32
rect 938 -38 950 -37
rect 938 -40 946 -38
rect 948 -40 950 -38
rect 938 -41 950 -40
rect 954 -38 960 -33
rect 954 -40 957 -38
rect 959 -40 960 -38
rect 954 -41 960 -40
rect 946 -45 950 -41
rect 946 -46 960 -45
rect 946 -48 950 -46
rect 952 -48 960 -46
rect 946 -49 960 -48
rect 969 -52 973 -23
rect 993 -22 997 -20
rect 993 -24 994 -22
rect 996 -24 997 -22
rect 993 -29 997 -24
rect 984 -30 997 -29
rect 984 -32 988 -30
rect 990 -32 997 -30
rect 984 -33 997 -32
rect 1001 -29 1005 -20
rect 1024 -21 1028 -12
rect 1024 -23 1026 -21
rect 1001 -30 1014 -29
rect 1001 -32 1010 -30
rect 1012 -32 1014 -30
rect 1001 -33 1014 -32
rect 992 -38 1004 -37
rect 992 -40 1000 -38
rect 1002 -40 1004 -38
rect 992 -41 1004 -40
rect 1008 -38 1014 -33
rect 1008 -40 1011 -38
rect 1013 -40 1014 -38
rect 1008 -41 1014 -40
rect 1000 -45 1004 -41
rect 1000 -46 1014 -45
rect 1000 -48 1002 -46
rect 1004 -48 1014 -46
rect 1000 -49 1014 -48
rect 1024 -52 1028 -23
rect 1048 -22 1052 -20
rect 1048 -24 1049 -22
rect 1051 -24 1052 -22
rect 1048 -29 1052 -24
rect 1039 -30 1052 -29
rect 1039 -32 1043 -30
rect 1045 -32 1052 -30
rect 1039 -33 1052 -32
rect 1056 -29 1060 -20
rect 1077 -21 1081 -12
rect 1077 -23 1079 -21
rect 1056 -30 1069 -29
rect 1056 -32 1065 -30
rect 1067 -32 1069 -30
rect 1056 -33 1069 -32
rect 1047 -38 1059 -37
rect 1047 -40 1055 -38
rect 1057 -40 1059 -38
rect 1047 -41 1059 -40
rect 1063 -38 1069 -33
rect 1063 -40 1066 -38
rect 1068 -40 1069 -38
rect 1063 -41 1069 -40
rect 1055 -45 1059 -41
rect 1055 -46 1069 -45
rect 1055 -48 1059 -46
rect 1061 -48 1069 -46
rect 1055 -49 1069 -48
rect 1077 -52 1081 -23
rect 1101 -22 1105 -20
rect 1101 -24 1102 -22
rect 1104 -24 1105 -22
rect 1101 -29 1105 -24
rect 1092 -30 1105 -29
rect 1092 -32 1096 -30
rect 1098 -32 1105 -30
rect 1092 -33 1105 -32
rect 1109 -29 1113 -20
rect 1109 -30 1122 -29
rect 1109 -32 1118 -30
rect 1120 -32 1122 -30
rect 1109 -33 1122 -32
rect 1100 -38 1112 -37
rect 1100 -40 1108 -38
rect 1110 -40 1112 -38
rect 1100 -41 1112 -40
rect 1116 -38 1122 -33
rect 1116 -40 1119 -38
rect 1121 -40 1122 -38
rect 1116 -41 1122 -40
rect 1108 -45 1112 -41
rect 1108 -46 1122 -45
rect 1108 -48 1111 -46
rect 1113 -48 1122 -46
rect 1108 -49 1122 -48
rect -156 -53 -144 -52
rect -156 -55 -154 -53
rect -152 -54 -144 -53
rect -152 -55 -151 -54
rect -156 -56 -151 -55
rect -149 -56 -144 -54
rect -104 -53 -92 -52
rect -104 -55 -102 -53
rect -100 -54 -92 -53
rect -100 -55 -99 -54
rect -104 -56 -99 -55
rect -97 -56 -92 -54
rect -52 -53 -40 -52
rect -52 -55 -50 -53
rect -48 -54 -40 -53
rect -48 -55 -47 -54
rect -52 -56 -47 -55
rect -45 -56 -40 -54
rect 0 -53 12 -52
rect 0 -55 2 -53
rect 4 -54 12 -53
rect 4 -55 5 -54
rect 0 -56 5 -55
rect 7 -56 12 -54
rect 52 -53 64 -52
rect 52 -55 54 -53
rect 56 -55 64 -53
rect -156 -58 -144 -56
rect -104 -58 -92 -56
rect -52 -58 -40 -56
rect 0 -58 12 -56
rect 52 -57 57 -55
rect 59 -57 64 -55
rect 105 -53 117 -52
rect 105 -55 107 -53
rect 109 -55 117 -53
rect 52 -58 64 -57
rect 105 -57 110 -55
rect 112 -57 117 -55
rect 162 -54 174 -52
rect 162 -56 171 -54
rect 173 -56 174 -54
rect 105 -58 117 -57
rect 162 -58 174 -56
rect 182 -54 194 -52
rect 182 -56 191 -54
rect 193 -56 194 -54
rect 182 -58 194 -56
rect 202 -54 214 -52
rect 202 -56 211 -54
rect 213 -56 214 -54
rect 202 -58 214 -56
rect 224 -54 236 -52
rect 224 -56 233 -54
rect 235 -56 236 -54
rect 224 -58 236 -56
rect 246 -54 258 -52
rect 246 -56 255 -54
rect 257 -56 258 -54
rect 246 -58 258 -56
rect 268 -54 280 -52
rect 268 -56 277 -54
rect 279 -56 280 -54
rect 268 -58 280 -56
rect 293 -53 305 -52
rect 293 -55 295 -53
rect 297 -55 305 -53
rect 293 -58 305 -55
rect 346 -53 358 -52
rect 346 -55 348 -53
rect 350 -55 358 -53
rect 346 -57 351 -55
rect 353 -57 358 -55
rect 398 -53 410 -52
rect 398 -55 400 -53
rect 402 -55 410 -53
rect 346 -58 358 -57
rect 398 -57 403 -55
rect 405 -57 410 -55
rect 450 -53 462 -52
rect 450 -55 452 -53
rect 454 -55 462 -53
rect 398 -58 410 -57
rect 450 -57 455 -55
rect 457 -57 462 -55
rect 502 -53 514 -52
rect 502 -55 504 -53
rect 506 -55 514 -53
rect 450 -58 462 -57
rect 502 -57 507 -55
rect 509 -57 514 -55
rect 557 -54 558 -52
rect 560 -54 569 -52
rect 557 -56 566 -54
rect 568 -56 569 -54
rect 502 -58 514 -57
rect 557 -58 569 -56
rect 578 -54 590 -52
rect 578 -56 580 -54
rect 582 -56 587 -54
rect 589 -56 590 -54
rect 578 -58 590 -56
rect 601 -53 613 -52
rect 601 -55 603 -53
rect 605 -55 613 -53
rect 601 -57 607 -55
rect 609 -57 613 -55
rect 654 -53 666 -52
rect 654 -55 656 -53
rect 658 -54 666 -53
rect 658 -55 659 -54
rect 654 -56 659 -55
rect 661 -56 666 -54
rect 706 -53 718 -52
rect 706 -55 708 -53
rect 710 -55 718 -53
rect 601 -58 613 -57
rect 654 -58 666 -56
rect 706 -57 711 -55
rect 713 -57 718 -55
rect 758 -53 770 -52
rect 758 -55 760 -53
rect 762 -55 770 -53
rect 706 -58 718 -57
rect 758 -57 763 -55
rect 765 -57 770 -55
rect 810 -53 822 -52
rect 810 -55 812 -53
rect 814 -55 822 -53
rect 758 -58 770 -57
rect 810 -57 816 -55
rect 818 -57 822 -55
rect 862 -53 874 -52
rect 862 -55 864 -53
rect 866 -55 874 -53
rect 810 -58 822 -57
rect 862 -57 867 -55
rect 869 -57 874 -55
rect 915 -53 927 -52
rect 915 -55 917 -53
rect 919 -55 927 -53
rect 862 -58 874 -57
rect 915 -57 920 -55
rect 922 -57 927 -55
rect 969 -53 981 -52
rect 969 -55 971 -53
rect 973 -55 981 -53
rect 915 -58 927 -57
rect 969 -57 974 -55
rect 976 -57 981 -55
rect 1024 -53 1036 -52
rect 1024 -55 1026 -53
rect 1028 -55 1036 -53
rect 969 -58 981 -57
rect 1024 -57 1030 -55
rect 1032 -57 1036 -55
rect 1077 -53 1089 -52
rect 1077 -55 1079 -53
rect 1081 -55 1089 -53
rect 1024 -58 1036 -57
rect 1077 -57 1086 -55
rect 1088 -57 1089 -55
rect 1077 -58 1089 -57
rect -158 -64 1133 -63
rect -158 -66 -143 -64
rect -141 -66 -133 -64
rect -131 -66 -123 -64
rect -121 -66 -91 -64
rect -89 -66 -81 -64
rect -79 -66 -71 -64
rect -69 -66 -39 -64
rect -37 -66 -29 -64
rect -27 -66 -19 -64
rect -17 -66 13 -64
rect 15 -66 23 -64
rect 25 -66 33 -64
rect 35 -66 65 -64
rect 67 -66 75 -64
rect 77 -66 85 -64
rect 87 -66 118 -64
rect 120 -66 128 -64
rect 130 -66 138 -64
rect 140 -66 164 -64
rect 166 -66 174 -64
rect 176 -66 184 -64
rect 186 -66 194 -64
rect 196 -66 204 -64
rect 206 -66 214 -64
rect 216 -66 226 -64
rect 228 -66 236 -64
rect 238 -66 248 -64
rect 250 -66 258 -64
rect 260 -66 270 -64
rect 272 -66 280 -64
rect 282 -66 306 -64
rect 308 -66 316 -64
rect 318 -66 326 -64
rect 328 -66 359 -64
rect 361 -66 369 -64
rect 371 -66 379 -64
rect 381 -66 411 -64
rect 413 -66 421 -64
rect 423 -66 431 -64
rect 433 -66 463 -64
rect 465 -66 473 -64
rect 475 -66 483 -64
rect 485 -66 515 -64
rect 517 -66 525 -64
rect 527 -66 535 -64
rect 537 -66 559 -64
rect 561 -66 569 -64
rect 571 -66 580 -64
rect 582 -66 590 -64
rect 592 -66 614 -64
rect 616 -66 624 -64
rect 626 -66 634 -64
rect 636 -66 667 -64
rect 669 -66 677 -64
rect 679 -66 687 -64
rect 689 -66 719 -64
rect 721 -66 729 -64
rect 731 -66 739 -64
rect 741 -66 771 -64
rect 773 -66 781 -64
rect 783 -66 791 -64
rect 793 -66 823 -64
rect 825 -66 833 -64
rect 835 -66 843 -64
rect 845 -66 875 -64
rect 877 -66 885 -64
rect 887 -66 895 -64
rect 897 -66 928 -64
rect 930 -66 938 -64
rect 940 -66 948 -64
rect 950 -66 982 -64
rect 984 -66 992 -64
rect 994 -66 1002 -64
rect 1004 -66 1037 -64
rect 1039 -66 1047 -64
rect 1049 -66 1057 -64
rect 1059 -65 1090 -64
rect 1059 -66 1078 -65
rect -158 -67 1078 -66
rect 1080 -66 1090 -65
rect 1092 -66 1100 -64
rect 1102 -66 1110 -64
rect 1112 -66 1133 -64
rect 1080 -67 1133 -66
rect -158 -71 1133 -67
<< alu2 >>
rect 89 358 101 359
rect 89 356 90 358
rect 92 356 98 358
rect 100 356 101 358
rect 89 355 101 356
rect 44 350 310 351
rect -277 348 -273 349
rect -277 346 -276 348
rect -274 346 -273 348
rect 44 348 45 350
rect 47 348 185 350
rect 187 348 310 350
rect 44 347 310 348
rect -277 344 -273 346
rect -277 342 -276 344
rect -274 342 -273 344
rect -277 341 -273 342
rect -124 343 -52 347
rect -124 334 -120 343
rect -124 332 -123 334
rect -121 332 -120 334
rect -124 331 -120 332
rect -56 335 -52 343
rect 44 339 48 347
rect 306 346 310 347
rect 357 347 587 351
rect 357 346 362 347
rect 306 342 362 346
rect 583 346 587 347
rect 634 347 863 351
rect 634 346 639 347
rect 583 342 639 346
rect 44 338 51 339
rect 44 336 48 338
rect 50 336 51 338
rect 44 335 51 336
rect 178 338 270 339
rect 178 336 267 338
rect 269 336 270 338
rect 178 335 270 336
rect 306 335 310 342
rect 455 338 547 339
rect 455 336 544 338
rect 546 336 547 338
rect 455 335 547 336
rect 583 335 587 342
rect 731 338 823 339
rect 731 336 820 338
rect 822 336 823 338
rect 731 335 823 336
rect 859 335 863 347
rect 1008 338 1100 339
rect 1008 336 1097 338
rect 1099 336 1100 338
rect 1008 335 1100 336
rect -56 334 -32 335
rect -56 332 -35 334
rect -33 332 -32 334
rect 178 334 182 335
rect -56 331 -32 332
rect 1 332 11 333
rect -267 330 -128 331
rect 1 330 2 332
rect 4 330 8 332
rect 10 330 11 332
rect 178 332 179 334
rect 181 332 182 334
rect 178 331 182 332
rect 306 334 318 335
rect 306 332 315 334
rect 317 332 318 334
rect 306 331 318 332
rect 455 334 459 335
rect 455 332 456 334
rect 458 332 459 334
rect 455 331 459 332
rect 583 334 595 335
rect 583 332 592 334
rect 594 332 595 334
rect 583 331 595 332
rect 731 334 735 335
rect 731 332 732 334
rect 734 332 735 334
rect 731 331 735 332
rect 859 334 871 335
rect 859 332 868 334
rect 870 332 871 334
rect 859 331 871 332
rect 1008 334 1012 335
rect 1008 332 1009 334
rect 1011 332 1012 334
rect 1008 331 1012 332
rect -267 328 -131 330
rect -129 328 -128 330
rect -267 327 -128 328
rect -115 329 -100 330
rect 1 329 11 330
rect 44 329 123 330
rect -115 327 -112 329
rect -110 327 -104 329
rect -102 327 -100 329
rect 44 327 120 329
rect 122 327 123 329
rect -266 322 -262 327
rect -115 326 -100 327
rect 39 326 123 327
rect 208 329 218 330
rect 208 327 209 329
rect 211 327 215 329
rect 217 327 218 329
rect 208 326 218 327
rect 346 329 400 330
rect 346 327 397 329
rect 399 327 400 329
rect 346 326 400 327
rect 485 329 495 330
rect 485 327 486 329
rect 488 327 492 329
rect 494 327 495 329
rect 485 326 495 327
rect 623 329 676 330
rect 623 327 673 329
rect 675 327 676 329
rect 623 326 676 327
rect 761 329 771 330
rect 761 327 762 329
rect 764 327 768 329
rect 770 327 771 329
rect 761 326 771 327
rect 899 329 953 330
rect 899 327 950 329
rect 952 327 953 329
rect 899 326 953 327
rect 1038 329 1048 330
rect 1038 327 1039 329
rect 1041 327 1045 329
rect 1047 327 1048 329
rect 1038 326 1048 327
rect 39 324 40 326
rect 42 324 48 326
rect 39 323 48 324
rect 346 324 347 326
rect 349 324 350 326
rect 346 323 350 324
rect 623 324 624 326
rect 626 324 627 326
rect 623 323 627 324
rect 899 324 900 326
rect 902 324 903 326
rect 899 323 903 324
rect -266 320 -265 322
rect -263 320 -262 322
rect -266 319 -262 320
rect -227 322 -179 323
rect -227 320 -226 322
rect -224 320 -182 322
rect -180 320 -179 322
rect -227 319 -179 320
rect -165 321 -154 322
rect -165 319 -164 321
rect -162 319 -157 321
rect -155 319 -154 321
rect -165 318 -154 319
rect -134 321 -31 322
rect -134 319 -133 321
rect -131 319 -35 321
rect -33 319 -31 321
rect -134 318 -31 319
rect 79 321 141 322
rect 79 319 80 321
rect 82 319 138 321
rect 140 319 141 321
rect 79 318 141 319
rect 168 321 271 322
rect 168 319 169 321
rect 171 319 267 321
rect 269 319 271 321
rect 168 318 271 319
rect 331 321 335 323
rect 331 319 332 321
rect 334 319 335 321
rect -4 317 0 318
rect -4 315 -3 317
rect -1 315 0 317
rect 298 317 306 318
rect -290 313 -271 315
rect -215 313 -89 314
rect -290 311 -274 313
rect -272 311 -271 313
rect -290 309 -271 311
rect -266 312 -262 313
rect -266 310 -265 312
rect -263 310 -262 312
rect -215 311 -214 313
rect -212 311 -92 313
rect -90 311 -89 313
rect -215 310 -89 311
rect -45 313 -41 314
rect -45 311 -44 313
rect -42 311 -41 313
rect -266 266 -262 310
rect -45 309 -41 311
rect -45 307 -44 309
rect -42 307 -41 309
rect -45 306 -41 307
rect -4 290 0 315
rect 43 315 59 316
rect -85 289 0 290
rect -85 287 -84 289
rect -82 287 0 289
rect -85 286 0 287
rect 15 312 19 314
rect 15 310 16 312
rect 18 310 19 312
rect 43 313 44 315
rect 46 313 56 315
rect 58 313 59 315
rect 298 315 299 317
rect 301 315 303 317
rect 305 315 306 317
rect 298 314 306 315
rect 43 311 59 313
rect 87 313 213 314
rect 87 311 88 313
rect 90 311 210 313
rect 212 311 213 313
rect 87 310 213 311
rect 15 281 19 310
rect 257 309 268 310
rect 257 307 258 309
rect 260 307 262 309
rect 264 307 268 309
rect 257 305 268 307
rect 209 292 218 293
rect 163 290 172 292
rect 163 288 164 290
rect 166 288 169 290
rect 171 288 172 290
rect 209 290 211 292
rect 213 290 215 292
rect 217 290 218 292
rect 209 289 218 290
rect 263 292 326 293
rect 263 290 264 292
rect 266 290 323 292
rect 325 290 326 292
rect 263 289 326 290
rect 163 287 172 288
rect -162 280 19 281
rect -162 278 -161 280
rect -159 279 318 280
rect -159 278 211 279
rect -162 277 211 278
rect 213 277 314 279
rect 316 277 318 279
rect 15 276 318 277
rect -69 266 -41 267
rect -266 264 -265 266
rect -263 264 -262 266
rect -282 245 -278 246
rect -282 243 -281 245
rect -279 243 -278 245
rect -282 239 -278 243
rect -282 237 -281 239
rect -279 237 -278 239
rect -282 234 -278 237
rect -282 188 -278 189
rect -282 186 -281 188
rect -279 186 -278 188
rect -282 180 -278 186
rect -282 178 -281 180
rect -279 178 -278 180
rect -282 172 -278 178
rect -266 177 -262 264
rect -215 265 -89 266
rect -215 263 -214 265
rect -212 263 -92 265
rect -90 263 -89 265
rect -215 262 -89 263
rect -69 264 -68 266
rect -66 265 -41 266
rect -66 264 -44 265
rect -69 263 -44 264
rect -42 263 -41 265
rect 55 266 59 276
rect 259 271 268 272
rect 259 269 260 271
rect 262 269 264 271
rect 266 269 268 271
rect 259 268 268 269
rect 55 264 56 266
rect 58 264 59 266
rect 55 263 59 264
rect 87 265 213 266
rect 87 263 88 265
rect 90 263 210 265
rect 212 263 213 265
rect -69 262 -41 263
rect 87 262 213 263
rect 217 263 270 264
rect 1 261 19 262
rect 1 259 2 261
rect 4 259 16 261
rect 18 259 19 261
rect 1 258 19 259
rect 217 261 267 263
rect 269 261 270 263
rect 217 260 270 261
rect 310 260 314 276
rect 217 258 221 260
rect -165 257 -154 258
rect -227 256 -179 257
rect -227 254 -226 256
rect -224 254 -182 256
rect -180 254 -179 256
rect -165 255 -164 257
rect -162 255 -161 257
rect -159 255 -154 257
rect -165 254 -154 255
rect -134 257 -31 258
rect -134 255 -133 257
rect -131 255 -35 257
rect -33 255 -31 257
rect -134 254 -31 255
rect 79 257 141 258
rect 79 255 80 257
rect 82 255 138 257
rect 140 255 141 257
rect 79 254 141 255
rect 168 257 221 258
rect 168 255 169 257
rect 171 255 221 257
rect 310 256 318 260
rect 168 254 221 255
rect -227 253 -179 254
rect 226 252 306 253
rect 226 250 227 252
rect 229 250 303 252
rect 305 250 306 252
rect -89 249 -81 250
rect -89 247 -88 249
rect -86 247 -84 249
rect -82 247 -81 249
rect -89 246 -81 247
rect -4 249 0 250
rect -4 247 -3 249
rect -1 247 0 249
rect -124 244 -120 245
rect -124 242 -123 244
rect -121 242 -120 244
rect -124 233 -120 242
rect -56 244 -32 245
rect -56 242 -35 244
rect -33 242 -32 244
rect -56 241 -32 242
rect -56 233 -52 241
rect -124 229 -52 233
rect -4 220 0 247
rect -91 218 0 220
rect -91 216 -90 218
rect -88 216 0 218
rect -91 215 0 216
rect 15 249 19 250
rect 15 247 16 249
rect 18 247 19 249
rect -164 208 -160 210
rect 15 208 19 247
rect 39 249 136 250
rect 226 249 306 250
rect 314 249 318 256
rect 39 247 40 249
rect 42 247 133 249
rect 135 247 136 249
rect 39 246 136 247
rect 314 247 315 249
rect 317 247 318 249
rect 314 246 318 247
rect 331 257 335 319
rect 354 321 418 322
rect 354 319 415 321
rect 417 319 418 321
rect 354 318 418 319
rect 445 321 548 322
rect 445 319 446 321
rect 448 319 544 321
rect 546 319 548 321
rect 445 318 548 319
rect 608 321 612 323
rect 608 319 609 321
rect 611 319 612 321
rect 354 293 358 318
rect 575 317 583 318
rect 575 315 576 317
rect 578 315 580 317
rect 582 315 583 317
rect 575 314 583 315
rect 364 313 490 314
rect 364 311 365 313
rect 367 311 487 313
rect 489 311 490 313
rect 364 310 490 311
rect 534 309 538 310
rect 534 307 535 309
rect 537 307 538 309
rect 534 305 538 307
rect 534 303 535 305
rect 537 303 538 305
rect 534 298 538 303
rect 341 292 358 293
rect 341 290 343 292
rect 345 290 358 292
rect 341 289 358 290
rect 486 292 495 293
rect 486 290 488 292
rect 490 290 492 292
rect 494 290 495 292
rect 486 289 495 290
rect 540 292 603 293
rect 540 290 541 292
rect 543 290 600 292
rect 602 290 603 292
rect 540 289 603 290
rect 347 279 595 280
rect 347 277 348 279
rect 350 277 591 279
rect 593 277 595 279
rect 347 276 595 277
rect 536 271 545 272
rect 536 269 537 271
rect 539 269 541 271
rect 543 269 545 271
rect 536 268 545 269
rect 364 265 490 266
rect 364 263 365 265
rect 367 263 487 265
rect 489 263 490 265
rect 364 262 490 263
rect 494 263 547 264
rect 494 261 544 263
rect 546 261 547 263
rect 494 260 547 261
rect 587 260 591 276
rect 494 258 498 260
rect 331 255 332 257
rect 334 255 335 257
rect 178 244 270 245
rect 178 242 179 244
rect 181 242 267 244
rect 269 242 270 244
rect 43 241 51 242
rect 178 241 270 242
rect 43 239 44 241
rect 46 239 48 241
rect 50 239 51 241
rect 43 238 51 239
rect 290 233 294 234
rect 290 231 291 233
rect 293 231 294 233
rect 88 218 103 219
rect 88 217 100 218
rect 88 215 89 217
rect 91 216 100 217
rect 102 216 103 218
rect 91 215 103 216
rect 88 214 103 215
rect -164 207 19 208
rect -164 205 -163 207
rect -161 206 267 207
rect -161 205 236 206
rect -164 204 236 205
rect 238 204 264 206
rect 266 204 267 206
rect -266 175 -265 177
rect -263 175 -262 177
rect -227 178 -179 179
rect -227 176 -226 178
rect -224 176 -182 178
rect -180 176 -179 178
rect -227 175 -179 176
rect -164 177 -160 204
rect 15 203 267 204
rect -124 192 -52 196
rect -124 190 -120 192
rect -124 188 -123 190
rect -121 188 -120 190
rect -124 187 -120 188
rect -56 191 -52 192
rect 47 194 51 203
rect 47 192 48 194
rect 50 192 51 194
rect 47 191 51 192
rect 178 194 270 195
rect 178 192 267 194
rect 269 192 270 194
rect 178 191 270 192
rect -56 190 -32 191
rect -56 188 -35 190
rect -33 188 -32 190
rect 178 190 182 191
rect -56 187 -32 188
rect 1 188 11 189
rect 1 186 2 188
rect 4 186 8 188
rect 10 186 11 188
rect 178 188 179 190
rect 181 188 182 190
rect 178 187 182 188
rect 290 186 294 231
rect 322 216 326 218
rect 322 214 323 216
rect 325 214 326 216
rect -91 185 -83 186
rect 1 185 11 186
rect 38 185 140 186
rect -91 183 -90 185
rect -88 183 -86 185
rect -84 183 -83 185
rect -91 182 -83 183
rect 38 183 40 185
rect 42 183 137 185
rect 139 183 140 185
rect 38 182 140 183
rect 226 185 294 186
rect 306 206 310 207
rect 306 204 307 206
rect 309 204 310 206
rect 306 190 310 204
rect 306 189 318 190
rect 306 187 315 189
rect 317 187 318 189
rect 306 185 318 187
rect 226 183 227 185
rect 229 183 294 185
rect 226 182 294 183
rect -164 175 -163 177
rect -161 175 -160 177
rect -266 122 -262 175
rect -164 174 -160 175
rect -134 177 -31 178
rect -134 175 -133 177
rect -131 175 -35 177
rect -33 175 -31 177
rect -134 174 -31 175
rect 79 177 142 178
rect 79 175 80 177
rect 82 175 139 177
rect 141 175 142 177
rect 79 174 142 175
rect 168 177 271 178
rect 322 177 326 214
rect 168 175 169 177
rect 171 175 267 177
rect 269 175 271 177
rect 168 174 271 175
rect -4 173 0 174
rect 298 173 306 174
rect -4 171 -3 173
rect -1 171 0 173
rect -215 169 -89 170
rect -215 167 -214 169
rect -212 167 -92 169
rect -90 167 -89 169
rect -215 166 -89 167
rect -45 167 -20 168
rect -45 165 -44 167
rect -42 165 -28 167
rect -26 165 -20 167
rect -45 164 -20 165
rect -4 146 0 171
rect 43 172 59 173
rect 43 170 44 172
rect 46 170 56 172
rect 58 170 59 172
rect 298 171 299 173
rect 301 171 303 173
rect 305 171 306 173
rect 298 170 306 171
rect 310 172 326 177
rect 331 177 335 255
rect 346 257 418 258
rect 346 256 415 257
rect 346 254 347 256
rect 349 255 415 256
rect 417 255 418 257
rect 349 254 418 255
rect 445 257 498 258
rect 445 255 446 257
rect 448 255 498 257
rect 587 256 595 260
rect 445 254 498 255
rect 346 253 361 254
rect 503 252 583 253
rect 503 250 504 252
rect 506 250 580 252
rect 582 250 583 252
rect 406 249 413 250
rect 503 249 583 250
rect 591 249 595 256
rect 406 247 410 249
rect 412 247 413 249
rect 406 246 413 247
rect 591 247 592 249
rect 594 247 595 249
rect 591 246 595 247
rect 608 257 612 319
rect 631 321 694 322
rect 631 319 691 321
rect 693 319 694 321
rect 631 318 694 319
rect 721 321 824 322
rect 721 319 722 321
rect 724 319 820 321
rect 822 319 824 321
rect 721 318 824 319
rect 884 321 888 323
rect 884 319 885 321
rect 887 319 888 321
rect 631 293 635 318
rect 851 317 859 318
rect 851 315 852 317
rect 854 315 856 317
rect 858 315 859 317
rect 851 314 859 315
rect 640 313 766 314
rect 640 311 641 313
rect 643 311 763 313
rect 765 311 766 313
rect 640 310 766 311
rect 790 310 814 311
rect 790 308 791 310
rect 793 308 811 310
rect 813 308 814 310
rect 790 306 814 308
rect 618 292 635 293
rect 618 290 620 292
rect 622 290 635 292
rect 618 289 635 290
rect 762 292 771 293
rect 762 290 764 292
rect 766 290 768 292
rect 770 290 771 292
rect 762 289 771 290
rect 816 292 879 293
rect 816 290 817 292
rect 819 290 876 292
rect 878 290 879 292
rect 816 289 879 290
rect 624 279 867 280
rect 624 277 625 279
rect 627 277 867 279
rect 624 276 867 277
rect 812 271 821 272
rect 812 269 813 271
rect 815 269 817 271
rect 819 269 821 271
rect 812 268 821 269
rect 640 265 766 266
rect 640 263 641 265
rect 643 263 763 265
rect 765 263 766 265
rect 640 262 766 263
rect 770 263 823 264
rect 770 261 820 263
rect 822 261 823 263
rect 770 260 823 261
rect 863 260 867 276
rect 770 258 774 260
rect 608 255 609 257
rect 611 255 612 257
rect 409 219 413 246
rect 455 244 547 245
rect 455 242 456 244
rect 458 242 544 244
rect 546 242 547 244
rect 455 241 547 242
rect 359 218 413 219
rect 340 216 413 218
rect 340 214 341 216
rect 343 214 413 216
rect 567 233 571 234
rect 567 231 568 233
rect 570 231 571 233
rect 340 212 361 214
rect 345 207 361 208
rect 345 205 347 207
rect 349 206 544 207
rect 349 205 541 206
rect 345 204 541 205
rect 543 204 544 206
rect 345 203 544 204
rect 455 194 547 195
rect 455 192 544 194
rect 546 192 547 194
rect 455 191 547 192
rect 455 190 459 191
rect 455 188 456 190
rect 458 188 459 190
rect 455 187 459 188
rect 567 186 571 231
rect 599 216 603 218
rect 599 214 600 216
rect 602 214 603 216
rect 346 185 417 186
rect 346 183 414 185
rect 416 183 417 185
rect 346 182 417 183
rect 503 185 571 186
rect 583 206 587 207
rect 583 204 584 206
rect 586 204 587 206
rect 583 190 587 204
rect 583 189 595 190
rect 583 187 592 189
rect 594 187 595 189
rect 583 185 595 187
rect 503 183 504 185
rect 506 183 571 185
rect 503 182 571 183
rect 346 180 347 182
rect 349 180 350 182
rect 346 179 350 180
rect 331 175 332 177
rect 334 175 335 177
rect 15 169 20 170
rect 43 169 59 170
rect 87 169 213 170
rect 15 167 16 169
rect 18 167 20 169
rect 15 165 20 167
rect 87 167 88 169
rect 90 167 210 169
rect 212 167 213 169
rect 87 166 213 167
rect -85 145 0 146
rect -85 143 -84 145
rect -82 143 0 145
rect -85 142 0 143
rect 16 136 20 165
rect 310 162 314 172
rect 257 161 314 162
rect 257 159 260 161
rect 262 159 314 161
rect 257 157 314 159
rect 331 167 335 175
rect 331 165 332 167
rect 334 165 335 167
rect 164 146 172 147
rect 164 144 165 146
rect 167 145 172 146
rect 167 144 169 145
rect 164 143 169 144
rect 171 143 172 145
rect 164 142 172 143
rect 263 144 327 145
rect 263 142 264 144
rect 266 142 324 144
rect 326 142 327 144
rect 263 141 327 142
rect -165 135 314 136
rect -165 134 253 135
rect -165 132 -164 134
rect -162 133 253 134
rect 255 133 311 135
rect 313 133 314 135
rect -162 132 314 133
rect -165 131 -50 132
rect -31 131 59 132
rect -45 127 -37 128
rect -45 126 -40 127
rect -45 124 -44 126
rect -42 125 -40 126
rect -38 125 -37 127
rect -42 124 -37 125
rect -45 123 -37 124
rect -266 120 -265 122
rect -263 120 -262 122
rect -282 92 -278 93
rect -282 90 -281 92
rect -279 90 -278 92
rect -282 89 -278 90
rect -282 87 -281 89
rect -279 87 -278 89
rect -282 86 -278 87
rect -283 53 -278 54
rect -283 51 -282 53
rect -280 51 -278 53
rect -283 50 -278 51
rect -283 48 -282 50
rect -280 48 -278 50
rect -283 47 -278 48
rect -266 33 -262 120
rect -215 121 -89 122
rect -41 121 -37 123
rect 54 121 59 131
rect 257 127 267 128
rect 257 125 260 127
rect 262 125 264 127
rect 266 125 267 127
rect 257 124 267 125
rect -215 119 -214 121
rect -212 119 -92 121
rect -90 119 -89 121
rect -215 118 -89 119
rect 54 119 56 121
rect 58 119 59 121
rect 1 117 19 118
rect 54 117 59 119
rect 87 121 213 122
rect 87 119 88 121
rect 90 119 210 121
rect 212 119 213 121
rect 87 118 213 119
rect 217 119 270 120
rect 217 117 267 119
rect 269 117 270 119
rect 1 115 2 117
rect 4 115 16 117
rect 18 115 19 117
rect 1 114 19 115
rect 217 116 270 117
rect 309 117 313 132
rect 217 114 221 116
rect -165 113 -154 114
rect -227 112 -179 113
rect -227 110 -226 112
rect -224 110 -182 112
rect -180 110 -179 112
rect -165 111 -164 113
rect -162 111 -157 113
rect -155 111 -154 113
rect -165 110 -154 111
rect -134 113 -31 114
rect -134 111 -133 113
rect -131 111 -35 113
rect -33 111 -31 113
rect -134 110 -31 111
rect 79 113 141 114
rect 79 111 80 113
rect 82 111 138 113
rect 140 111 141 113
rect 79 110 141 111
rect 168 113 221 114
rect 309 113 318 117
rect 168 111 169 113
rect 171 111 221 113
rect 168 110 221 111
rect -227 109 -179 110
rect 226 108 306 109
rect 226 106 227 108
rect 229 106 303 108
rect 305 106 306 108
rect -89 105 -81 106
rect -89 103 -88 105
rect -86 103 -84 105
rect -82 103 -81 105
rect -89 102 -81 103
rect -4 105 0 106
rect -4 103 -3 105
rect -1 103 0 105
rect -124 100 -120 101
rect -124 98 -123 100
rect -121 98 -120 100
rect -124 89 -120 98
rect -56 100 -32 101
rect -56 98 -35 100
rect -33 98 -32 100
rect -56 97 -32 98
rect -56 89 -52 97
rect -124 85 -52 89
rect -4 73 0 103
rect -85 72 0 73
rect -85 70 -84 72
rect -82 70 0 72
rect -85 68 0 70
rect 16 105 20 106
rect 16 103 17 105
rect 19 103 20 105
rect 16 63 20 103
rect 39 105 135 106
rect 226 105 306 106
rect 314 105 318 113
rect 39 103 40 105
rect 42 103 131 105
rect 133 103 135 105
rect 39 102 135 103
rect 314 103 315 105
rect 317 103 318 105
rect 314 102 318 103
rect 331 113 335 165
rect 355 177 419 178
rect 355 175 416 177
rect 418 175 419 177
rect 355 174 419 175
rect 445 177 548 178
rect 599 177 603 214
rect 445 175 446 177
rect 448 175 544 177
rect 546 175 548 177
rect 445 174 548 175
rect 355 145 359 174
rect 575 173 583 174
rect 575 171 576 173
rect 578 171 580 173
rect 582 171 583 173
rect 575 170 583 171
rect 587 172 603 177
rect 608 177 612 255
rect 623 257 694 258
rect 623 256 691 257
rect 623 254 624 256
rect 626 255 691 256
rect 693 255 694 257
rect 626 254 694 255
rect 721 257 774 258
rect 721 255 722 257
rect 724 255 774 257
rect 863 256 871 260
rect 721 254 774 255
rect 623 253 638 254
rect 779 252 859 253
rect 779 250 780 252
rect 782 250 856 252
rect 858 250 859 252
rect 684 249 689 250
rect 779 249 859 250
rect 867 249 871 256
rect 684 247 686 249
rect 688 247 689 249
rect 684 246 689 247
rect 867 247 868 249
rect 870 247 871 249
rect 867 246 871 247
rect 884 257 888 319
rect 907 321 971 322
rect 907 319 968 321
rect 970 319 971 321
rect 907 318 971 319
rect 998 321 1101 322
rect 998 319 999 321
rect 1001 319 1097 321
rect 1099 319 1101 321
rect 998 318 1101 319
rect 907 293 911 318
rect 1128 317 1136 318
rect 1128 315 1129 317
rect 1131 315 1133 317
rect 1135 315 1136 317
rect 1128 314 1136 315
rect 917 313 1043 314
rect 917 311 918 313
rect 920 311 1040 313
rect 1042 311 1043 313
rect 917 310 1043 311
rect 1087 308 1091 309
rect 1087 306 1088 308
rect 1090 306 1091 308
rect 1087 299 1091 306
rect 1087 297 1088 299
rect 1090 297 1091 299
rect 894 292 911 293
rect 894 290 896 292
rect 898 290 911 292
rect 894 289 911 290
rect 1039 292 1048 293
rect 1039 290 1041 292
rect 1043 290 1045 292
rect 1047 290 1048 292
rect 1039 289 1048 290
rect 1087 286 1091 297
rect 1082 274 1093 275
rect 1082 272 1084 274
rect 1086 272 1090 274
rect 1092 272 1093 274
rect 1082 270 1093 272
rect 917 265 1043 266
rect 917 263 918 265
rect 920 263 1040 265
rect 1042 263 1043 265
rect 917 262 1043 263
rect 1047 263 1100 264
rect 1047 261 1097 263
rect 1099 261 1100 263
rect 1047 260 1100 261
rect 1047 258 1051 260
rect 884 255 885 257
rect 887 255 888 257
rect 685 218 689 246
rect 731 244 823 245
rect 731 242 732 244
rect 734 242 820 244
rect 822 242 823 244
rect 731 241 823 242
rect 617 216 689 218
rect 617 214 618 216
rect 620 214 689 216
rect 617 212 689 214
rect 843 233 847 234
rect 843 231 844 233
rect 846 231 847 233
rect 622 207 638 208
rect 622 205 624 207
rect 626 206 820 207
rect 626 205 817 206
rect 622 204 817 205
rect 819 204 820 206
rect 622 203 820 204
rect 731 194 823 195
rect 731 192 820 194
rect 822 192 823 194
rect 731 191 823 192
rect 731 190 735 191
rect 731 188 732 190
rect 734 188 735 190
rect 731 187 735 188
rect 843 186 847 231
rect 875 216 879 218
rect 875 214 876 216
rect 878 214 879 216
rect 623 185 693 186
rect 623 183 690 185
rect 692 183 693 185
rect 623 182 693 183
rect 779 185 847 186
rect 859 206 863 207
rect 859 204 860 206
rect 862 204 863 206
rect 859 190 863 204
rect 859 189 871 190
rect 859 187 868 189
rect 870 187 871 189
rect 859 185 871 187
rect 779 183 780 185
rect 782 183 847 185
rect 779 182 847 183
rect 623 180 624 182
rect 626 180 627 182
rect 623 179 627 180
rect 608 175 609 177
rect 611 175 612 177
rect 364 169 490 170
rect 364 167 365 169
rect 367 167 487 169
rect 489 167 490 169
rect 364 166 490 167
rect 587 162 591 172
rect 534 161 591 162
rect 534 159 537 161
rect 539 159 591 161
rect 534 157 591 159
rect 339 144 359 145
rect 339 142 340 144
rect 342 142 359 144
rect 339 141 359 142
rect 540 144 604 145
rect 540 142 541 144
rect 543 142 601 144
rect 603 142 604 144
rect 540 141 604 142
rect 346 135 591 136
rect 346 133 347 135
rect 349 133 588 135
rect 590 133 591 135
rect 346 132 591 133
rect 534 127 544 128
rect 534 125 537 127
rect 539 125 541 127
rect 543 125 544 127
rect 534 124 544 125
rect 364 121 490 122
rect 364 119 365 121
rect 367 119 487 121
rect 489 119 490 121
rect 364 118 490 119
rect 494 119 547 120
rect 494 117 544 119
rect 546 117 547 119
rect 494 116 547 117
rect 586 117 590 132
rect 494 114 498 116
rect 331 111 332 113
rect 334 111 335 113
rect 178 100 270 101
rect 178 98 179 100
rect 181 98 267 100
rect 269 98 270 100
rect 43 97 51 98
rect 178 97 270 98
rect 43 95 44 97
rect 46 95 48 97
rect 50 95 51 97
rect 43 94 51 95
rect 289 89 293 90
rect 289 87 290 89
rect 292 87 293 89
rect 88 73 102 74
rect 88 71 89 73
rect 91 71 99 73
rect 101 71 102 73
rect 88 70 102 71
rect -164 62 20 63
rect -164 60 -163 62
rect -161 60 20 62
rect -164 59 20 60
rect -266 31 -265 33
rect -263 31 -262 33
rect -227 34 -179 35
rect -227 32 -226 34
rect -224 32 -182 34
rect -180 32 -179 34
rect -227 31 -179 32
rect -164 33 -160 59
rect -124 49 -52 55
rect -124 46 -120 49
rect -124 44 -123 46
rect -121 44 -120 46
rect -124 43 -120 44
rect -56 47 -52 49
rect 16 51 20 59
rect 53 63 265 64
rect 53 61 261 63
rect 263 61 265 63
rect 53 60 265 61
rect 53 51 57 60
rect 16 50 57 51
rect 16 48 48 50
rect 50 48 57 50
rect 16 47 57 48
rect 178 50 270 51
rect 178 48 267 50
rect 269 48 270 50
rect 178 47 270 48
rect -56 46 -32 47
rect -56 44 -35 46
rect -33 44 -32 46
rect 178 46 182 47
rect -56 43 -32 44
rect 1 44 11 45
rect 1 42 2 44
rect 4 42 8 44
rect 10 42 11 44
rect 178 44 179 46
rect 181 44 182 46
rect 178 43 182 44
rect 289 42 293 87
rect 322 72 326 73
rect 322 70 323 72
rect 325 70 326 72
rect 306 63 310 64
rect 306 61 307 63
rect 309 61 310 63
rect 306 50 310 61
rect 306 49 318 50
rect 306 47 315 49
rect 317 47 318 49
rect 306 46 318 47
rect -89 41 -81 42
rect 1 41 11 42
rect 128 41 136 42
rect -89 39 -88 41
rect -86 39 -84 41
rect -82 39 -81 41
rect -89 38 -81 39
rect 128 39 129 41
rect 131 39 133 41
rect 135 39 136 41
rect 128 38 136 39
rect 225 41 294 42
rect 225 39 226 41
rect 228 39 294 41
rect 225 38 294 39
rect 322 36 326 70
rect -164 31 -163 33
rect -161 31 -160 33
rect -266 29 -262 31
rect -164 30 -160 31
rect -134 33 -31 34
rect 79 33 141 34
rect -134 31 -133 33
rect -131 31 -35 33
rect -33 31 -31 33
rect -134 30 -31 31
rect -5 31 0 33
rect -5 29 -3 31
rect -1 29 0 31
rect 79 31 80 33
rect 82 31 138 33
rect 140 31 141 33
rect 79 30 141 31
rect 168 33 271 34
rect 168 31 169 33
rect 171 31 193 33
rect 195 31 267 33
rect 269 31 271 33
rect 168 30 271 31
rect 298 33 306 34
rect 298 31 299 33
rect 301 31 303 33
rect 305 31 306 33
rect 298 30 306 31
rect 310 31 326 36
rect 331 33 335 111
rect 350 113 418 114
rect 350 111 415 113
rect 417 111 418 113
rect 350 110 418 111
rect 445 113 498 114
rect 586 113 595 117
rect 445 111 446 113
rect 448 111 498 113
rect 445 110 498 111
rect 346 109 354 110
rect 346 107 347 109
rect 349 107 354 109
rect 346 106 354 107
rect 503 108 583 109
rect 503 106 504 108
rect 506 106 580 108
rect 582 106 583 108
rect 407 105 412 106
rect 503 105 583 106
rect 591 105 595 113
rect 407 103 408 105
rect 410 103 412 105
rect 407 74 412 103
rect 591 103 592 105
rect 594 103 595 105
rect 591 102 595 103
rect 608 113 612 175
rect 632 177 695 178
rect 632 175 692 177
rect 694 175 695 177
rect 632 174 695 175
rect 721 177 824 178
rect 875 177 879 214
rect 721 175 722 177
rect 724 175 820 177
rect 822 175 824 177
rect 721 174 824 175
rect 632 145 636 174
rect 851 173 859 174
rect 851 171 852 173
rect 854 171 856 173
rect 858 171 859 173
rect 851 170 859 171
rect 863 172 879 177
rect 884 177 888 255
rect 899 257 971 258
rect 899 256 968 257
rect 899 254 900 256
rect 902 255 968 256
rect 970 255 971 257
rect 902 254 971 255
rect 998 257 1051 258
rect 998 255 999 257
rect 1001 255 1051 257
rect 998 254 1051 255
rect 899 253 914 254
rect 1056 252 1136 253
rect 1056 250 1057 252
rect 1059 250 1133 252
rect 1135 250 1136 252
rect 959 249 966 250
rect 1056 249 1136 250
rect 959 247 963 249
rect 965 247 966 249
rect 959 246 966 247
rect 962 219 966 246
rect 1008 244 1100 245
rect 1008 242 1009 244
rect 1011 242 1097 244
rect 1099 242 1100 244
rect 1008 241 1100 242
rect 912 218 966 219
rect 893 216 966 218
rect 893 214 894 216
rect 896 214 966 216
rect 1120 233 1124 234
rect 1120 231 1121 233
rect 1123 231 1124 233
rect 893 212 914 214
rect 1008 194 1100 195
rect 1008 192 1097 194
rect 1099 192 1100 194
rect 1008 191 1100 192
rect 1008 190 1012 191
rect 1008 188 1009 190
rect 1011 188 1012 190
rect 1008 187 1012 188
rect 1120 186 1124 231
rect 899 185 970 186
rect 899 183 967 185
rect 969 183 970 185
rect 899 182 970 183
rect 1056 185 1124 186
rect 1056 183 1057 185
rect 1059 183 1124 185
rect 1056 182 1124 183
rect 899 180 900 182
rect 902 180 903 182
rect 899 179 903 180
rect 884 175 885 177
rect 887 175 888 177
rect 640 169 766 170
rect 640 167 641 169
rect 643 167 763 169
rect 765 167 766 169
rect 640 166 766 167
rect 863 162 867 172
rect 810 161 867 162
rect 810 159 813 161
rect 815 159 867 161
rect 810 157 867 159
rect 616 144 636 145
rect 616 142 617 144
rect 619 142 636 144
rect 616 141 636 142
rect 816 144 880 145
rect 816 142 817 144
rect 819 142 877 144
rect 879 142 880 144
rect 816 141 880 142
rect 623 135 867 136
rect 623 133 624 135
rect 626 133 864 135
rect 866 133 867 135
rect 623 132 867 133
rect 810 127 820 128
rect 810 125 813 127
rect 815 125 817 127
rect 819 125 820 127
rect 810 124 820 125
rect 640 121 766 122
rect 640 119 641 121
rect 643 119 763 121
rect 765 119 766 121
rect 640 118 766 119
rect 770 119 823 120
rect 770 117 820 119
rect 822 117 823 119
rect 770 116 823 117
rect 862 117 866 132
rect 770 114 774 116
rect 608 111 609 113
rect 611 111 612 113
rect 455 100 547 101
rect 455 98 456 100
rect 458 98 544 100
rect 546 98 547 100
rect 455 97 547 98
rect 350 73 412 74
rect 339 72 412 73
rect 339 70 340 72
rect 342 70 412 72
rect 566 89 570 90
rect 566 87 567 89
rect 569 87 570 89
rect 339 69 354 70
rect 339 64 352 65
rect 339 62 345 64
rect 347 63 542 64
rect 347 62 538 63
rect 339 61 538 62
rect 540 61 542 63
rect 348 60 542 61
rect 455 50 547 51
rect 455 48 544 50
rect 546 48 547 50
rect 455 47 547 48
rect 455 46 459 47
rect 455 44 456 46
rect 458 44 459 46
rect 455 43 459 44
rect 566 42 570 87
rect 608 88 612 111
rect 634 113 694 114
rect 634 111 691 113
rect 693 111 694 113
rect 634 110 694 111
rect 721 113 774 114
rect 862 113 871 117
rect 721 111 722 113
rect 724 111 774 113
rect 721 110 774 111
rect 623 109 638 110
rect 623 107 624 109
rect 626 107 638 109
rect 623 106 638 107
rect 779 108 859 109
rect 779 106 780 108
rect 782 106 856 108
rect 858 106 859 108
rect 681 105 688 106
rect 779 105 859 106
rect 867 105 871 113
rect 681 103 684 105
rect 686 103 688 105
rect 681 102 688 103
rect 867 103 868 105
rect 870 103 871 105
rect 867 102 871 103
rect 884 113 888 175
rect 908 177 972 178
rect 908 175 969 177
rect 971 175 972 177
rect 908 174 972 175
rect 998 177 1101 178
rect 998 175 999 177
rect 1001 175 1097 177
rect 1099 175 1101 177
rect 998 174 1101 175
rect 908 145 912 174
rect 1128 173 1136 174
rect 1128 171 1129 173
rect 1131 171 1133 173
rect 1135 171 1136 173
rect 1128 170 1136 171
rect 917 169 1043 170
rect 917 167 918 169
rect 920 167 1040 169
rect 1042 167 1043 169
rect 917 166 1043 167
rect 1087 164 1091 166
rect 1087 162 1088 164
rect 1090 162 1091 164
rect 1087 146 1091 162
rect 892 144 912 145
rect 892 142 893 144
rect 895 142 912 144
rect 892 141 912 142
rect 939 145 1091 146
rect 939 143 940 145
rect 942 143 1091 145
rect 939 141 1091 143
rect 1083 129 1093 131
rect 1083 127 1084 129
rect 1086 127 1090 129
rect 1092 127 1093 129
rect 1083 125 1093 127
rect 917 121 1043 122
rect 917 119 918 121
rect 920 119 1040 121
rect 1042 119 1043 121
rect 917 118 1043 119
rect 1047 119 1100 120
rect 1047 117 1097 119
rect 1099 117 1100 119
rect 1047 116 1100 117
rect 1047 114 1051 116
rect 884 111 885 113
rect 887 111 888 113
rect 608 86 609 88
rect 611 86 612 88
rect 599 72 603 73
rect 599 70 600 72
rect 602 70 603 72
rect 583 63 587 64
rect 583 61 584 63
rect 586 61 587 63
rect 583 50 587 61
rect 583 49 595 50
rect 583 47 592 49
rect 594 47 595 49
rect 583 46 595 47
rect 346 41 413 42
rect 346 39 410 41
rect 412 39 413 41
rect 346 37 347 39
rect 349 38 413 39
rect 502 41 571 42
rect 502 39 503 41
rect 505 39 571 41
rect 502 38 571 39
rect 349 37 350 38
rect 346 36 350 37
rect 599 36 603 70
rect 331 31 332 33
rect 334 31 335 33
rect -5 26 0 29
rect 43 27 59 28
rect -215 25 -89 26
rect -215 23 -214 25
rect -212 23 -92 25
rect -90 23 -89 25
rect -215 22 -89 23
rect -45 22 -10 24
rect -45 20 -44 22
rect -42 20 -13 22
rect -11 20 -10 22
rect -45 19 -10 20
rect -80 0 -65 1
rect -132 -2 -128 0
rect -132 -4 -131 -2
rect -129 -4 -128 -2
rect -132 -21 -128 -4
rect -132 -23 -131 -21
rect -129 -23 -128 -21
rect -132 -25 -128 -23
rect -80 -2 -68 0
rect -66 -2 -65 0
rect -80 -3 -65 -2
rect -80 -21 -76 -3
rect -5 -6 -1 26
rect 43 25 44 27
rect 46 25 56 27
rect 58 25 59 27
rect 14 24 22 25
rect 14 22 15 24
rect 17 22 19 24
rect 21 22 22 24
rect 43 23 59 25
rect 87 25 213 26
rect 87 23 88 25
rect 90 23 210 25
rect 212 23 213 25
rect 87 22 213 23
rect 257 23 261 24
rect 14 21 22 22
rect 257 21 258 23
rect 260 21 261 23
rect 257 20 261 21
rect 310 20 314 31
rect 331 30 335 31
rect 355 33 418 34
rect 355 31 357 33
rect 359 31 415 33
rect 417 31 418 33
rect 355 30 418 31
rect 445 33 548 34
rect 445 31 446 33
rect 448 31 544 33
rect 546 31 548 33
rect 445 30 548 31
rect 575 33 583 34
rect 575 31 576 33
rect 578 31 580 33
rect 582 31 583 33
rect 575 30 583 31
rect 587 31 603 36
rect 608 33 612 86
rect 683 73 687 102
rect 731 100 823 101
rect 731 98 732 100
rect 734 98 820 100
rect 822 98 823 100
rect 731 97 823 98
rect 616 72 687 73
rect 616 70 617 72
rect 619 70 687 72
rect 616 69 687 70
rect 842 89 846 90
rect 842 87 843 89
rect 845 87 846 89
rect 616 64 641 65
rect 616 62 622 64
rect 624 63 818 64
rect 624 62 814 63
rect 616 61 814 62
rect 816 61 818 63
rect 637 60 818 61
rect 731 50 823 51
rect 731 48 820 50
rect 822 48 823 50
rect 731 47 823 48
rect 731 46 735 47
rect 731 44 732 46
rect 734 44 735 46
rect 731 43 735 44
rect 842 42 846 87
rect 875 72 879 73
rect 875 70 876 72
rect 878 70 879 72
rect 859 63 863 64
rect 859 61 860 63
rect 862 61 863 63
rect 859 50 863 61
rect 859 49 871 50
rect 859 47 868 49
rect 870 47 871 49
rect 859 46 871 47
rect 623 41 689 42
rect 623 39 686 41
rect 688 39 689 41
rect 623 37 624 39
rect 626 38 689 39
rect 778 41 847 42
rect 778 39 779 41
rect 781 39 847 41
rect 778 38 847 39
rect 626 37 627 38
rect 623 36 627 37
rect 875 36 879 70
rect 608 31 609 33
rect 611 31 612 33
rect 364 25 490 26
rect 364 23 365 25
rect 367 23 487 25
rect 489 23 490 25
rect 364 22 490 23
rect 534 23 538 24
rect 31 18 43 19
rect 31 17 35 18
rect 31 15 32 17
rect 34 16 35 17
rect 37 16 43 18
rect 257 16 314 20
rect 534 21 535 23
rect 537 21 538 23
rect 534 20 538 21
rect 587 20 591 31
rect 608 30 612 31
rect 632 33 694 34
rect 632 31 634 33
rect 636 31 691 33
rect 693 31 694 33
rect 632 30 694 31
rect 721 33 824 34
rect 721 31 722 33
rect 724 31 820 33
rect 822 31 824 33
rect 721 30 824 31
rect 851 33 859 34
rect 851 31 852 33
rect 854 31 856 33
rect 858 31 859 33
rect 851 30 859 31
rect 863 31 879 36
rect 884 46 888 111
rect 903 113 971 114
rect 903 111 968 113
rect 970 111 971 113
rect 903 110 971 111
rect 998 113 1051 114
rect 998 111 999 113
rect 1001 111 1051 113
rect 998 110 1051 111
rect 899 109 907 110
rect 899 107 900 109
rect 902 107 907 109
rect 899 106 907 107
rect 1056 108 1136 109
rect 1056 106 1057 108
rect 1059 106 1133 108
rect 1135 106 1136 108
rect 960 105 965 106
rect 1056 105 1136 106
rect 960 103 961 105
rect 963 103 965 105
rect 960 74 965 103
rect 1008 100 1100 101
rect 1008 98 1009 100
rect 1011 98 1097 100
rect 1099 98 1100 100
rect 1008 97 1100 98
rect 1119 89 1123 90
rect 1119 87 1120 89
rect 1122 87 1123 89
rect 903 73 965 74
rect 892 72 965 73
rect 892 70 893 72
rect 895 70 965 72
rect 1067 74 1080 75
rect 1067 72 1069 74
rect 1071 72 1080 74
rect 1067 70 1074 72
rect 1076 70 1080 72
rect 892 69 907 70
rect 1067 69 1080 70
rect 884 44 885 46
rect 887 44 888 46
rect 884 33 888 44
rect 1008 50 1100 51
rect 1008 48 1097 50
rect 1099 48 1100 50
rect 1008 47 1100 48
rect 1008 46 1012 47
rect 1008 44 1009 46
rect 1011 44 1012 46
rect 1008 43 1012 44
rect 1119 42 1123 87
rect 899 41 966 42
rect 899 39 963 41
rect 965 39 966 41
rect 899 37 900 39
rect 902 38 966 39
rect 1055 41 1124 42
rect 1055 39 1056 41
rect 1058 39 1124 41
rect 1055 38 1124 39
rect 902 37 903 38
rect 899 36 903 37
rect 884 31 885 33
rect 887 31 888 33
rect 640 25 766 26
rect 640 23 641 25
rect 643 23 763 25
rect 765 23 766 25
rect 640 22 766 23
rect 810 23 814 24
rect 534 16 591 20
rect 810 21 811 23
rect 813 21 814 23
rect 810 20 814 21
rect 863 20 867 31
rect 884 30 888 31
rect 908 33 971 34
rect 908 31 910 33
rect 912 31 968 33
rect 970 31 971 33
rect 908 30 971 31
rect 998 33 1101 34
rect 998 31 999 33
rect 1001 31 1097 33
rect 1099 31 1101 33
rect 998 30 1101 31
rect 1128 30 1132 32
rect 1128 28 1129 30
rect 1131 28 1132 30
rect 917 25 1043 26
rect 917 23 918 25
rect 920 23 1040 25
rect 1042 23 1043 25
rect 917 22 1043 23
rect 810 16 867 20
rect 1087 20 1091 21
rect 1087 18 1088 20
rect 1090 18 1091 20
rect 34 15 43 16
rect 31 13 43 15
rect 163 5 172 7
rect 1087 5 1091 18
rect 1128 7 1132 28
rect 128 4 138 5
rect 128 2 129 4
rect 131 2 134 4
rect 136 2 138 4
rect 128 1 138 2
rect 163 3 164 5
rect 166 3 169 5
rect 171 3 172 5
rect 163 1 172 3
rect 671 4 682 5
rect 671 2 672 4
rect 674 2 682 4
rect 671 1 682 2
rect -5 -10 133 -6
rect -80 -23 -79 -21
rect -77 -23 -76 -21
rect -80 -24 -76 -23
rect -28 -15 -24 -14
rect -28 -17 -27 -15
rect -25 -17 -24 -15
rect -28 -21 -24 -17
rect -28 -23 -27 -21
rect -25 -23 -24 -21
rect 76 -22 80 -20
rect -28 -25 -24 -23
rect 24 -23 28 -22
rect 24 -25 25 -23
rect 27 -25 28 -23
rect 24 -29 28 -25
rect 24 -31 25 -29
rect 27 -31 28 -29
rect 76 -24 77 -22
rect 79 -24 80 -22
rect 76 -27 80 -24
rect 129 -22 133 -10
rect 625 -15 629 -6
rect 625 -17 626 -15
rect 628 -17 629 -15
rect 129 -24 130 -22
rect 132 -24 133 -22
rect 129 -25 133 -24
rect 183 -22 321 -20
rect 183 -24 318 -22
rect 320 -24 321 -22
rect 625 -23 629 -17
rect 76 -29 77 -27
rect 79 -29 80 -27
rect 183 -26 184 -24
rect 186 -25 321 -24
rect 186 -26 188 -25
rect 526 -26 530 -24
rect 625 -25 626 -23
rect 628 -25 629 -23
rect 678 -21 682 1
rect 790 2 794 5
rect 790 0 791 2
rect 793 0 794 2
rect 1048 1 1091 5
rect 1101 2 1132 7
rect 730 -3 734 -1
rect 724 -4 734 -3
rect 724 -6 725 -4
rect 727 -6 734 -4
rect 724 -8 734 -6
rect 678 -23 679 -21
rect 681 -23 682 -21
rect 678 -25 682 -23
rect 730 -22 734 -8
rect 790 -11 794 0
rect 730 -24 731 -22
rect 733 -24 734 -22
rect 730 -25 734 -24
rect 782 -15 794 -11
rect 886 -3 890 0
rect 886 -5 887 -3
rect 889 -5 890 -3
rect 782 -22 786 -15
rect 782 -24 783 -22
rect 785 -24 786 -22
rect 782 -25 786 -24
rect 834 -16 845 -15
rect 834 -18 841 -16
rect 843 -18 845 -16
rect 834 -20 845 -18
rect 834 -22 838 -20
rect 834 -24 835 -22
rect 837 -24 838 -22
rect 834 -25 838 -24
rect 886 -22 890 -5
rect 1018 -4 1022 -2
rect 1018 -6 1019 -4
rect 1021 -6 1022 -4
rect 886 -24 887 -22
rect 889 -24 890 -22
rect 625 -26 629 -25
rect 183 -28 188 -26
rect 422 -27 426 -26
rect 422 -29 423 -27
rect 425 -29 426 -27
rect 526 -28 527 -26
rect 529 -28 530 -26
rect 886 -27 890 -24
rect 939 -17 943 -15
rect 939 -19 940 -17
rect 942 -19 943 -17
rect 939 -22 943 -19
rect 1018 -20 1022 -6
rect 939 -24 940 -22
rect 942 -24 943 -22
rect 939 -26 943 -24
rect 993 -22 1022 -20
rect 993 -24 994 -22
rect 996 -24 1022 -22
rect 993 -25 1022 -24
rect 1048 -22 1052 1
rect 1048 -24 1049 -22
rect 1051 -24 1052 -22
rect 1048 -25 1052 -24
rect 1101 -22 1105 2
rect 1101 -24 1102 -22
rect 1104 -24 1105 -22
rect 1101 -25 1105 -24
rect 76 -31 80 -29
rect 204 -30 208 -29
rect 204 -31 213 -30
rect 24 -32 28 -31
rect 204 -33 205 -31
rect 207 -33 210 -31
rect 212 -33 213 -31
rect 204 -34 213 -33
rect 229 -31 236 -30
rect 229 -33 230 -31
rect 232 -33 233 -31
rect 235 -33 236 -31
rect 229 -34 236 -33
rect 248 -31 306 -29
rect 248 -33 250 -31
rect 252 -33 299 -31
rect 301 -33 306 -31
rect 361 -30 371 -29
rect 361 -32 362 -30
rect 364 -32 368 -30
rect 370 -32 371 -30
rect 248 -34 306 -33
rect 332 -35 338 -32
rect 361 -33 371 -32
rect 420 -30 426 -29
rect 420 -32 421 -30
rect 423 -32 426 -30
rect 420 -33 426 -32
rect 465 -30 476 -29
rect 465 -32 466 -30
rect 468 -32 473 -30
rect 475 -32 476 -30
rect 465 -33 476 -32
rect 526 -30 530 -28
rect 526 -32 527 -30
rect 529 -32 530 -30
rect 526 -33 530 -32
rect -158 -38 166 -37
rect -158 -40 -114 -38
rect -112 -40 -62 -38
rect -60 -40 -10 -38
rect -8 -40 42 -38
rect 44 -40 94 -38
rect 96 -40 147 -38
rect 149 -40 166 -38
rect -158 -41 166 -40
rect 162 -45 166 -41
rect -158 -46 155 -45
rect -158 -48 -120 -46
rect -118 -48 -69 -46
rect -67 -48 -16 -46
rect -14 -48 35 -46
rect 37 -48 87 -46
rect 89 -48 140 -46
rect 142 -48 155 -46
rect -158 -49 155 -48
rect -152 -54 -148 -53
rect -152 -56 -151 -54
rect -149 -56 -148 -54
rect -152 -80 -148 -56
rect -100 -54 -96 -53
rect -100 -56 -99 -54
rect -97 -56 -96 -54
rect -100 -83 -96 -56
rect -48 -54 -44 -53
rect -48 -56 -47 -54
rect -45 -56 -44 -54
rect -48 -79 -44 -56
rect 4 -54 8 -53
rect 4 -56 5 -54
rect 7 -56 8 -54
rect 4 -82 8 -56
rect 55 -55 60 -53
rect 55 -57 57 -55
rect 59 -57 60 -55
rect 55 -83 60 -57
rect 109 -55 114 -54
rect 109 -57 110 -55
rect 112 -57 114 -55
rect 109 -83 114 -57
rect 151 -68 155 -49
rect 162 -47 163 -45
rect 165 -47 166 -45
rect 170 -38 174 -35
rect 332 -37 335 -35
rect 337 -37 338 -35
rect 565 -36 569 -34
rect 332 -38 547 -37
rect 170 -40 171 -38
rect 173 -40 174 -38
rect 170 -43 174 -40
rect 276 -39 287 -38
rect 276 -41 277 -39
rect 279 -41 284 -39
rect 286 -41 287 -39
rect 276 -42 287 -41
rect 293 -40 304 -39
rect 293 -42 294 -40
rect 296 -42 298 -40
rect 300 -42 304 -40
rect 332 -40 335 -38
rect 337 -40 388 -38
rect 390 -40 440 -38
rect 442 -40 492 -38
rect 494 -40 544 -38
rect 546 -40 547 -38
rect 332 -41 547 -40
rect 565 -38 566 -36
rect 568 -38 569 -36
rect 202 -43 206 -42
rect 293 -43 304 -42
rect 170 -45 171 -43
rect 173 -45 174 -43
rect 170 -47 174 -45
rect 182 -45 191 -43
rect 182 -47 183 -45
rect 185 -47 188 -45
rect 190 -47 191 -45
rect 162 -51 166 -47
rect 182 -49 191 -47
rect 202 -45 203 -43
rect 205 -45 206 -43
rect 246 -45 250 -44
rect 202 -47 206 -45
rect 202 -49 203 -47
rect 205 -49 206 -47
rect 202 -50 206 -49
rect 224 -46 237 -45
rect 224 -48 225 -46
rect 227 -47 237 -46
rect 227 -48 234 -47
rect 224 -49 234 -48
rect 236 -49 237 -47
rect 224 -50 237 -49
rect 246 -47 247 -45
rect 249 -47 250 -45
rect 246 -48 250 -47
rect 246 -50 247 -48
rect 249 -50 250 -48
rect 246 -51 250 -50
rect 268 -46 272 -43
rect 268 -48 269 -46
rect 271 -48 272 -46
rect 268 -49 272 -48
rect 268 -51 269 -49
rect 271 -51 272 -49
rect 293 -51 297 -43
rect 565 -45 569 -38
rect 586 -38 1131 -37
rect 586 -40 587 -38
rect 589 -40 643 -38
rect 645 -40 696 -38
rect 698 -40 748 -38
rect 750 -40 800 -38
rect 802 -40 852 -38
rect 854 -40 904 -38
rect 906 -40 957 -38
rect 959 -40 1011 -38
rect 1013 -40 1066 -38
rect 1068 -40 1119 -38
rect 1121 -40 1131 -38
rect 586 -41 1131 -40
rect 328 -46 540 -45
rect 328 -48 329 -46
rect 331 -48 382 -46
rect 384 -48 433 -46
rect 435 -48 486 -46
rect 488 -48 537 -46
rect 539 -48 540 -46
rect 565 -46 1131 -45
rect 565 -48 643 -46
rect 645 -48 690 -46
rect 692 -48 741 -46
rect 743 -48 794 -46
rect 796 -48 845 -46
rect 847 -48 897 -46
rect 899 -48 950 -46
rect 952 -48 1002 -46
rect 1004 -48 1059 -46
rect 1061 -48 1111 -46
rect 1113 -48 1131 -46
rect 328 -49 540 -48
rect 162 -53 163 -51
rect 165 -53 166 -51
rect 268 -52 272 -51
rect 162 -54 166 -53
rect 328 -68 332 -49
rect 151 -73 332 -68
rect 350 -55 354 -54
rect 350 -57 351 -55
rect 353 -57 354 -55
rect 350 -81 354 -57
rect 402 -55 406 -54
rect 402 -57 403 -55
rect 405 -57 406 -55
rect 402 -80 406 -57
rect 454 -55 458 -54
rect 454 -57 455 -55
rect 457 -57 458 -55
rect 454 -80 458 -57
rect 506 -55 510 -54
rect 506 -57 507 -55
rect 509 -57 510 -55
rect 506 -81 510 -57
rect 536 -68 540 -49
rect 557 -49 561 -48
rect 565 -49 1131 -48
rect 557 -51 558 -49
rect 560 -51 561 -49
rect 557 -52 561 -51
rect 557 -54 558 -52
rect 560 -54 561 -52
rect 557 -57 561 -54
rect 578 -54 583 -53
rect 657 -54 662 -53
rect 578 -56 580 -54
rect 582 -56 583 -54
rect 578 -68 583 -56
rect 536 -73 583 -68
rect 606 -55 610 -54
rect 606 -57 607 -55
rect 609 -57 610 -55
rect 606 -81 610 -57
rect 657 -56 659 -54
rect 661 -56 662 -54
rect 657 -79 662 -56
rect 709 -55 714 -54
rect 709 -57 711 -55
rect 713 -57 714 -55
rect 709 -83 714 -57
rect 762 -55 766 -54
rect 762 -57 763 -55
rect 765 -57 766 -55
rect 762 -79 766 -57
rect 814 -55 819 -54
rect 814 -57 816 -55
rect 818 -57 819 -55
rect 814 -84 819 -57
rect 865 -55 870 -54
rect 865 -57 867 -55
rect 869 -57 870 -55
rect 865 -84 870 -57
rect 918 -55 923 -54
rect 918 -57 920 -55
rect 922 -57 923 -55
rect 918 -81 923 -57
rect 973 -55 977 -54
rect 973 -57 974 -55
rect 976 -57 977 -55
rect 973 -81 977 -57
rect 1028 -55 1033 -54
rect 1028 -57 1030 -55
rect 1032 -57 1033 -55
rect 1028 -81 1033 -57
rect 1085 -55 1089 -54
rect 1085 -57 1086 -55
rect 1088 -57 1089 -55
rect 1073 -65 1081 -63
rect 1073 -67 1074 -65
rect 1076 -67 1078 -65
rect 1080 -67 1081 -65
rect 1073 -69 1081 -67
rect 1085 -81 1089 -57
<< alu3 >>
rect 84 358 93 359
rect 84 357 90 358
rect 84 355 85 357
rect 87 356 90 357
rect 92 356 93 358
rect 87 355 93 356
rect 84 354 93 355
rect 29 350 48 351
rect -277 348 5 349
rect -277 346 -276 348
rect -274 346 5 348
rect 29 348 31 350
rect 33 348 45 350
rect 47 348 48 350
rect 29 347 48 348
rect 184 350 192 351
rect 184 348 185 350
rect 187 348 188 350
rect 190 348 192 350
rect 184 347 192 348
rect -277 345 5 346
rect -165 339 -161 340
rect -165 337 -164 339
rect -162 337 -161 339
rect -165 322 -161 337
rect 1 332 5 345
rect -133 330 -124 331
rect 1 330 2 332
rect 4 330 5 332
rect -133 328 -131 330
rect -129 329 -109 330
rect -129 328 -112 329
rect -133 327 -112 328
rect -110 327 -109 329
rect -128 326 -109 327
rect -290 321 -161 322
rect -290 319 -164 321
rect -162 319 -161 321
rect -290 318 -161 319
rect -290 317 -162 318
rect -52 316 -41 317
rect -52 314 -51 316
rect -49 314 -41 316
rect -52 313 -41 314
rect -52 312 -44 313
rect -45 311 -44 312
rect -42 311 -41 313
rect -45 310 -41 311
rect -85 289 -81 290
rect -85 287 -84 289
rect -82 287 -81 289
rect -288 280 -158 283
rect -288 279 -161 280
rect -162 278 -161 279
rect -159 278 -158 280
rect -282 273 -278 274
rect -282 271 -281 273
rect -279 271 -278 273
rect -282 245 -278 271
rect -162 257 -158 278
rect -162 255 -161 257
rect -159 255 -158 257
rect -162 254 -158 255
rect -85 249 -81 287
rect -61 273 -3 274
rect -61 271 -60 273
rect -58 271 -6 273
rect -4 271 -3 273
rect -61 270 -3 271
rect -85 247 -84 249
rect -82 247 -81 249
rect -85 246 -81 247
rect -69 266 -65 267
rect -69 264 -68 266
rect -66 264 -65 266
rect -282 243 -281 245
rect -279 243 -278 245
rect -282 241 -278 243
rect -91 218 -87 220
rect -91 216 -90 218
rect -88 216 -87 218
rect -286 207 -160 210
rect -286 205 -163 207
rect -161 205 -160 207
rect -286 203 -160 205
rect -91 185 -87 216
rect -91 183 -90 185
rect -88 183 -87 185
rect -91 182 -87 183
rect -282 180 -278 181
rect -282 178 -281 180
rect -279 178 -278 180
rect -282 175 -278 178
rect -282 173 -281 175
rect -279 173 -278 175
rect -282 164 -278 173
rect -85 145 -81 146
rect -85 143 -84 145
rect -82 143 -81 145
rect -287 134 -161 136
rect -287 132 -164 134
rect -162 132 -161 134
rect -165 113 -161 132
rect -165 111 -164 113
rect -162 111 -161 113
rect -165 110 -161 111
rect -85 105 -81 143
rect -85 103 -84 105
rect -82 103 -81 105
rect -85 102 -81 103
rect -282 89 -274 90
rect -282 87 -281 89
rect -279 87 -277 89
rect -275 87 -274 89
rect -282 86 -274 87
rect -85 72 -81 73
rect -85 70 -84 72
rect -82 70 -81 72
rect -290 62 -160 63
rect -290 60 -163 62
rect -161 60 -160 62
rect -290 59 -160 60
rect -283 50 -278 51
rect -283 48 -282 50
rect -280 48 -278 50
rect -283 46 -278 48
rect -283 44 -282 46
rect -280 44 -278 46
rect -283 43 -278 44
rect -85 41 -81 70
rect -85 39 -84 41
rect -82 39 -81 41
rect -85 38 -81 39
rect -69 0 -65 264
rect 1 261 5 330
rect 214 329 218 330
rect 214 327 215 329
rect 217 327 218 329
rect 1 259 2 261
rect 4 259 5 261
rect 1 188 5 259
rect 1 186 2 188
rect 4 186 5 188
rect -29 167 -20 168
rect -29 165 -28 167
rect -26 165 -24 167
rect -22 165 -20 167
rect -29 164 -20 165
rect -41 127 -37 128
rect -41 125 -40 127
rect -38 125 -37 127
rect -41 123 -37 125
rect -41 121 -40 123
rect -38 121 -37 123
rect -41 120 -37 121
rect 1 117 5 186
rect 1 115 2 117
rect 4 115 5 117
rect 1 44 5 115
rect 1 42 2 44
rect 4 42 5 44
rect 1 41 5 42
rect 43 315 47 316
rect 43 313 44 315
rect 46 313 47 315
rect 43 273 47 313
rect 214 292 218 327
rect 491 329 495 330
rect 491 327 492 329
rect 494 327 495 329
rect 302 317 306 318
rect 302 315 303 317
rect 305 315 306 317
rect 257 309 268 310
rect 257 307 262 309
rect 264 307 265 309
rect 267 307 268 309
rect 257 305 268 307
rect 167 291 177 292
rect 167 290 174 291
rect 167 288 169 290
rect 171 289 174 290
rect 176 289 177 291
rect 214 290 215 292
rect 217 290 218 292
rect 214 289 218 290
rect 263 292 267 293
rect 263 290 264 292
rect 266 290 267 292
rect 171 288 177 289
rect 167 287 177 288
rect 43 271 44 273
rect 46 271 47 273
rect 43 241 47 271
rect 43 239 44 241
rect 46 239 47 241
rect 43 172 47 239
rect 210 279 214 280
rect 210 277 211 279
rect 213 277 214 279
rect 84 217 92 219
rect 84 215 85 217
rect 87 215 89 217
rect 91 215 92 217
rect 84 214 92 215
rect 43 170 44 172
rect 46 170 47 172
rect 43 97 47 170
rect 168 145 177 147
rect 168 143 169 145
rect 171 143 173 145
rect 175 143 177 145
rect 168 142 177 143
rect 43 95 44 97
rect 46 95 47 97
rect 43 27 47 95
rect 84 73 92 74
rect 84 71 85 73
rect 87 71 89 73
rect 91 71 92 73
rect 84 70 92 71
rect 43 25 44 27
rect 46 25 47 27
rect 18 24 28 25
rect -132 -2 -99 0
rect -132 -4 -131 -2
rect -129 -4 -102 -2
rect -100 -4 -99 -2
rect -69 -2 -68 0
rect -66 -2 -65 0
rect -69 -3 -65 -2
rect -14 22 -10 24
rect -14 20 -13 22
rect -11 20 -10 22
rect 18 22 19 24
rect 21 22 24 24
rect 26 22 28 24
rect 43 23 47 25
rect 128 41 132 42
rect 128 39 129 41
rect 131 39 132 41
rect 18 21 28 22
rect -14 -2 -10 20
rect 34 18 43 19
rect 34 16 35 18
rect 37 16 39 18
rect 41 16 43 18
rect 34 14 43 16
rect 128 4 132 39
rect 158 33 200 34
rect 158 31 160 33
rect 162 31 193 33
rect 195 32 200 33
rect 195 31 197 32
rect 158 30 197 31
rect 199 30 200 32
rect 158 29 200 30
rect 128 2 129 4
rect 131 2 132 4
rect 128 1 132 2
rect 167 5 177 7
rect 167 3 169 5
rect 171 3 174 5
rect 176 3 177 5
rect 167 1 177 3
rect 210 4 214 277
rect 263 271 267 290
rect 263 269 264 271
rect 266 269 267 271
rect 263 268 267 269
rect 302 252 306 315
rect 322 292 346 293
rect 491 292 495 327
rect 767 329 771 330
rect 767 327 768 329
rect 770 327 771 329
rect 579 317 583 318
rect 579 315 580 317
rect 582 315 583 317
rect 534 305 538 310
rect 534 303 535 305
rect 537 303 538 305
rect 534 302 538 303
rect 534 300 535 302
rect 537 300 538 302
rect 534 298 538 300
rect 322 290 323 292
rect 325 290 343 292
rect 345 290 346 292
rect 410 290 414 292
rect 322 289 346 290
rect 409 288 411 290
rect 413 288 414 290
rect 491 290 492 292
rect 494 290 495 292
rect 491 289 495 290
rect 540 292 544 293
rect 540 290 541 292
rect 543 290 544 292
rect 312 279 353 280
rect 312 277 314 279
rect 316 277 348 279
rect 350 277 353 279
rect 312 276 353 277
rect 312 275 325 276
rect 302 250 303 252
rect 305 250 306 252
rect 302 249 306 250
rect 322 216 344 218
rect 322 214 323 216
rect 325 214 341 216
rect 343 214 344 216
rect 322 212 344 214
rect 210 2 211 4
rect 213 2 214 4
rect 187 -2 191 0
rect 210 -1 214 2
rect 235 206 240 209
rect 345 207 350 208
rect 235 204 236 206
rect 238 204 240 206
rect 235 2 240 204
rect 263 206 347 207
rect 263 204 264 206
rect 266 204 307 206
rect 309 205 347 206
rect 349 205 350 207
rect 309 204 350 205
rect 263 203 350 204
rect 302 173 306 174
rect 302 171 303 173
rect 305 171 306 173
rect 263 144 267 145
rect 263 142 264 144
rect 266 142 267 144
rect 235 0 237 2
rect 239 0 240 2
rect 235 -1 240 0
rect 252 135 256 136
rect 252 133 253 135
rect 255 133 256 135
rect 252 3 256 133
rect 263 127 267 142
rect 263 125 264 127
rect 266 125 267 127
rect 263 124 267 125
rect 302 108 306 171
rect 328 167 335 168
rect 328 165 329 167
rect 331 165 332 167
rect 334 165 335 167
rect 328 162 335 165
rect 323 144 343 145
rect 323 142 324 144
rect 326 142 340 144
rect 342 142 343 144
rect 323 141 343 142
rect 310 135 352 136
rect 310 133 311 135
rect 313 133 347 135
rect 349 133 352 135
rect 310 132 352 133
rect 302 106 303 108
rect 305 106 306 108
rect 302 105 306 106
rect 409 75 414 288
rect 540 271 544 290
rect 540 269 541 271
rect 543 269 544 271
rect 540 268 544 269
rect 579 252 583 315
rect 599 292 623 293
rect 599 290 600 292
rect 602 290 620 292
rect 622 290 623 292
rect 599 289 623 290
rect 767 292 771 327
rect 1044 329 1048 330
rect 1044 327 1045 329
rect 1047 327 1048 329
rect 855 317 859 318
rect 855 315 856 317
rect 858 315 859 317
rect 767 290 768 292
rect 770 290 771 292
rect 767 289 771 290
rect 790 310 794 311
rect 790 308 791 310
rect 793 308 794 310
rect 724 288 729 289
rect 724 286 726 288
rect 728 286 729 288
rect 589 279 630 280
rect 589 277 591 279
rect 593 277 625 279
rect 627 277 630 279
rect 589 276 630 277
rect 589 275 602 276
rect 579 250 580 252
rect 582 250 583 252
rect 579 249 583 250
rect 599 216 621 218
rect 599 214 600 216
rect 602 214 618 216
rect 620 214 621 216
rect 599 212 621 214
rect 622 207 627 208
rect 540 206 624 207
rect 540 204 541 206
rect 543 204 584 206
rect 586 205 624 206
rect 626 205 627 207
rect 586 204 627 205
rect 540 203 627 204
rect 579 173 583 174
rect 579 171 580 173
rect 582 171 583 173
rect 540 144 544 145
rect 540 142 541 144
rect 543 142 544 144
rect 540 127 544 142
rect 540 125 541 127
rect 543 125 544 127
rect 540 124 544 125
rect 579 108 583 171
rect 600 144 620 145
rect 600 142 601 144
rect 603 142 617 144
rect 619 142 620 144
rect 600 141 620 142
rect 587 135 629 136
rect 587 133 588 135
rect 590 133 624 135
rect 626 133 629 135
rect 587 132 629 133
rect 579 106 580 108
rect 582 106 583 108
rect 579 105 583 106
rect 593 89 612 90
rect 593 87 603 89
rect 605 88 612 89
rect 605 87 609 88
rect 593 86 609 87
rect 611 86 612 88
rect 593 85 612 86
rect 322 72 343 73
rect 322 70 323 72
rect 325 70 340 72
rect 342 70 343 72
rect 322 69 343 70
rect 409 72 554 75
rect 671 73 675 75
rect 409 70 550 72
rect 552 70 554 72
rect 409 68 554 70
rect 599 72 620 73
rect 599 70 600 72
rect 602 70 617 72
rect 619 70 620 72
rect 599 69 620 70
rect 671 71 672 73
rect 674 71 675 73
rect 308 64 348 65
rect 585 64 625 65
rect 260 63 345 64
rect 260 61 261 63
rect 263 61 270 63
rect 272 61 307 63
rect 309 62 345 63
rect 347 62 348 64
rect 309 61 348 62
rect 260 60 348 61
rect 536 63 622 64
rect 536 61 538 63
rect 540 61 584 63
rect 586 62 622 63
rect 624 62 625 64
rect 586 61 625 62
rect 536 60 625 61
rect 302 33 306 34
rect 302 31 303 33
rect 305 31 306 33
rect 302 30 306 31
rect 354 33 361 34
rect 354 31 357 33
rect 359 31 361 33
rect 354 30 361 31
rect 579 33 583 34
rect 579 31 580 33
rect 582 31 583 33
rect 579 30 583 31
rect 631 33 638 34
rect 631 31 634 33
rect 636 31 638 33
rect 631 30 638 31
rect 302 26 358 30
rect 579 26 635 30
rect 252 1 253 3
rect 255 1 256 3
rect 671 4 675 71
rect 671 2 672 4
rect 674 2 675 4
rect 671 1 675 2
rect 252 -1 256 1
rect -132 -5 -99 -4
rect -14 -6 80 -2
rect -28 -15 -20 -14
rect -28 -17 -27 -15
rect -25 -17 -23 -15
rect -21 -17 -20 -15
rect -28 -18 -20 -17
rect 24 -17 28 -16
rect 24 -19 25 -17
rect 27 -19 28 -17
rect 24 -23 28 -19
rect 24 -25 25 -23
rect 27 -25 28 -23
rect 24 -26 28 -25
rect 76 -22 80 -6
rect 76 -24 77 -22
rect 79 -24 80 -22
rect 76 -26 80 -24
rect 187 -4 188 -2
rect 190 -4 191 -2
rect 170 -43 174 -41
rect 170 -45 171 -43
rect 173 -45 174 -43
rect 162 -51 166 -48
rect 162 -53 163 -51
rect 165 -53 166 -51
rect 162 -59 166 -53
rect 162 -61 163 -59
rect 165 -61 166 -59
rect 162 -63 166 -61
rect 170 -61 174 -45
rect 187 -45 191 -4
rect 724 -4 729 286
rect 790 2 794 308
rect 816 292 820 293
rect 816 290 817 292
rect 819 290 820 292
rect 816 271 820 290
rect 816 269 817 271
rect 819 269 820 271
rect 816 268 820 269
rect 855 252 859 315
rect 875 292 899 293
rect 875 290 876 292
rect 878 290 896 292
rect 898 290 899 292
rect 875 289 899 290
rect 1044 292 1048 327
rect 1132 317 1136 318
rect 1132 315 1133 317
rect 1135 315 1136 317
rect 1044 290 1045 292
rect 1047 290 1048 292
rect 1044 289 1048 290
rect 1087 299 1091 309
rect 1087 297 1088 299
rect 1090 297 1091 299
rect 1087 289 1091 297
rect 1087 287 1088 289
rect 1090 287 1091 289
rect 1087 286 1091 287
rect 855 250 856 252
rect 858 250 859 252
rect 855 249 859 250
rect 927 274 1093 275
rect 927 272 1084 274
rect 1086 272 1093 274
rect 927 271 1093 272
rect 875 216 897 218
rect 875 214 876 216
rect 878 214 894 216
rect 896 214 897 216
rect 875 212 897 214
rect 816 206 863 207
rect 816 204 817 206
rect 819 204 860 206
rect 862 204 863 206
rect 816 203 863 204
rect 855 173 859 174
rect 855 171 856 173
rect 858 171 859 173
rect 816 144 820 145
rect 816 142 817 144
rect 819 142 820 144
rect 816 127 820 142
rect 816 125 817 127
rect 819 125 820 127
rect 816 124 820 125
rect 855 108 859 171
rect 876 144 896 145
rect 876 142 877 144
rect 879 142 893 144
rect 895 142 896 144
rect 876 141 896 142
rect 863 135 867 136
rect 863 133 864 135
rect 866 133 867 135
rect 863 132 867 133
rect 855 106 856 108
rect 858 106 859 108
rect 855 105 859 106
rect 875 72 896 73
rect 875 70 876 72
rect 878 70 893 72
rect 895 70 896 72
rect 875 69 896 70
rect 812 63 863 64
rect 812 61 814 63
rect 816 61 860 63
rect 862 61 863 63
rect 812 60 863 61
rect 868 46 888 47
rect 868 44 876 46
rect 878 44 885 46
rect 887 44 888 46
rect 868 43 888 44
rect 855 33 859 34
rect 855 31 856 33
rect 858 31 859 33
rect 855 30 859 31
rect 907 33 914 34
rect 907 31 910 33
rect 912 31 914 33
rect 907 30 914 31
rect 855 26 911 30
rect 790 0 791 2
rect 793 0 794 2
rect 790 -2 794 0
rect 840 3 845 5
rect 840 1 842 3
rect 844 1 845 3
rect 724 -6 725 -4
rect 727 -6 729 -4
rect 625 -7 629 -6
rect 204 -13 365 -8
rect 515 -10 530 -8
rect 515 -12 517 -10
rect 519 -12 530 -10
rect 515 -13 530 -12
rect 204 -31 208 -13
rect 232 -22 352 -20
rect 232 -24 347 -22
rect 349 -24 352 -22
rect 232 -25 352 -24
rect 232 -30 236 -25
rect 204 -33 205 -31
rect 207 -33 208 -31
rect 204 -34 208 -33
rect 229 -31 236 -30
rect 229 -33 233 -31
rect 235 -33 236 -31
rect 229 -34 236 -33
rect 298 -31 330 -29
rect 298 -33 299 -31
rect 301 -33 327 -31
rect 329 -33 330 -31
rect 361 -30 365 -13
rect 370 -22 423 -20
rect 370 -24 371 -22
rect 373 -24 423 -22
rect 370 -25 423 -24
rect 361 -32 362 -30
rect 364 -32 365 -30
rect 361 -33 365 -32
rect 419 -29 423 -25
rect 419 -30 424 -29
rect 419 -32 421 -30
rect 423 -32 424 -30
rect 298 -34 330 -33
rect 419 -34 424 -32
rect 456 -30 469 -29
rect 456 -31 466 -30
rect 456 -33 458 -31
rect 460 -32 466 -31
rect 468 -32 469 -30
rect 460 -33 469 -32
rect 526 -30 530 -13
rect 625 -9 626 -7
rect 628 -9 629 -7
rect 724 -8 729 -6
rect 625 -15 629 -9
rect 625 -17 626 -15
rect 628 -17 629 -15
rect 625 -26 629 -17
rect 840 -16 845 1
rect 927 0 931 271
rect 1082 270 1093 271
rect 1132 252 1136 315
rect 1132 250 1133 252
rect 1135 250 1136 252
rect 1132 249 1136 250
rect 1132 173 1136 174
rect 1132 171 1133 173
rect 1135 171 1136 173
rect 886 -3 931 0
rect 886 -5 887 -3
rect 889 -5 931 -3
rect 886 -6 931 -5
rect 939 145 943 148
rect 939 143 940 145
rect 942 143 943 145
rect 840 -18 841 -16
rect 843 -18 845 -16
rect 840 -20 845 -18
rect 939 -17 943 143
rect 1018 131 1023 132
rect 1018 129 1093 131
rect 1018 127 1084 129
rect 1086 127 1093 129
rect 1018 125 1093 127
rect 1018 68 1023 125
rect 1132 108 1136 171
rect 1132 106 1133 108
rect 1135 106 1136 108
rect 1132 105 1136 106
rect 1073 72 1077 74
rect 1073 70 1074 72
rect 1076 70 1077 72
rect 1018 -4 1022 68
rect 1018 -6 1019 -4
rect 1021 -6 1022 -4
rect 1018 -7 1022 -6
rect 939 -19 940 -17
rect 942 -19 943 -17
rect 939 -26 943 -19
rect 526 -32 527 -30
rect 529 -32 530 -30
rect 526 -33 530 -32
rect 456 -34 469 -33
rect 334 -35 338 -34
rect 268 -39 274 -36
rect 334 -37 335 -35
rect 337 -37 338 -35
rect 268 -41 271 -39
rect 273 -41 274 -39
rect 187 -47 188 -45
rect 190 -47 191 -45
rect 202 -43 214 -42
rect 202 -45 203 -43
rect 205 -45 211 -43
rect 213 -45 214 -43
rect 246 -45 256 -44
rect 202 -47 214 -45
rect 233 -46 241 -45
rect 233 -47 238 -46
rect 187 -49 191 -47
rect 233 -49 234 -47
rect 236 -48 238 -47
rect 240 -48 241 -46
rect 246 -47 247 -45
rect 249 -47 253 -45
rect 255 -47 256 -45
rect 246 -48 256 -47
rect 268 -46 274 -41
rect 282 -39 293 -38
rect 282 -41 284 -39
rect 286 -41 289 -39
rect 291 -41 293 -39
rect 282 -43 293 -41
rect 297 -40 304 -39
rect 297 -42 298 -40
rect 300 -42 301 -40
rect 303 -42 304 -40
rect 297 -43 304 -42
rect 334 -41 338 -37
rect 334 -43 335 -41
rect 337 -43 338 -41
rect 334 -44 338 -43
rect 268 -48 269 -46
rect 271 -48 274 -46
rect 236 -49 241 -48
rect 268 -49 274 -48
rect 557 -49 561 -48
rect 233 -50 241 -49
rect 557 -50 558 -49
rect 283 -51 558 -50
rect 560 -51 561 -49
rect 283 -52 561 -51
rect 283 -54 285 -52
rect 287 -54 561 -52
rect 283 -55 334 -54
rect 347 -55 561 -54
rect 170 -62 338 -61
rect 170 -64 335 -62
rect 337 -64 338 -62
rect 170 -65 338 -64
rect 1073 -65 1077 70
rect 1073 -67 1074 -65
rect 1076 -67 1077 -65
rect 1073 -72 1077 -67
<< alu4 >>
rect 84 357 88 358
rect 84 355 85 357
rect 87 355 88 357
rect -165 350 39 351
rect -165 348 31 350
rect 33 348 39 350
rect -165 347 39 348
rect -165 339 -161 347
rect -165 337 -164 339
rect -162 337 -161 339
rect -165 333 -161 337
rect -52 316 -48 317
rect -52 314 -51 316
rect -49 314 -48 316
rect -282 273 -57 274
rect -282 271 -281 273
rect -279 271 -60 273
rect -58 271 -57 273
rect -282 270 -57 271
rect -282 175 -278 181
rect -282 173 -281 175
rect -279 173 -278 175
rect -282 167 -278 173
rect -282 165 -281 167
rect -279 165 -278 167
rect -282 164 -278 165
rect -278 89 -271 90
rect -278 87 -277 89
rect -275 87 -274 89
rect -272 87 -271 89
rect -278 86 -271 87
rect -283 46 -270 47
rect -283 44 -282 46
rect -280 44 -274 46
rect -272 44 -270 46
rect -283 43 -270 44
rect -52 1 -48 314
rect 29 278 34 347
rect -7 273 20 274
rect -7 271 -6 273
rect -4 271 17 273
rect 19 271 20 273
rect -7 270 20 271
rect 29 266 33 278
rect 37 273 47 274
rect 37 271 38 273
rect 40 271 44 273
rect 46 271 47 273
rect 37 270 47 271
rect -28 167 -20 168
rect -28 165 -24 167
rect -22 165 -20 167
rect -28 164 -20 165
rect -41 123 -37 124
rect -41 121 -40 123
rect -38 121 -37 123
rect -41 70 -37 121
rect -53 0 -48 1
rect -103 -2 -48 0
rect -42 1 -37 70
rect -42 -1 -40 1
rect -38 -1 -37 1
rect -42 -2 -37 -1
rect -103 -4 -102 -2
rect -100 -3 -48 -2
rect -100 -4 -49 -3
rect -103 -5 -49 -4
rect -24 -15 -20 164
rect 29 25 34 266
rect 84 217 88 355
rect 187 350 191 351
rect 187 348 188 350
rect 190 348 191 350
rect 84 215 85 217
rect 87 215 88 217
rect 84 73 88 215
rect 84 71 85 73
rect 87 71 88 73
rect 84 70 88 71
rect 172 291 177 292
rect 172 289 174 291
rect 176 289 177 291
rect 172 145 177 289
rect 172 143 173 145
rect 175 143 177 145
rect 21 24 34 25
rect 21 22 24 24
rect 26 22 34 24
rect 21 21 34 22
rect 39 33 164 34
rect 39 31 160 33
rect 162 31 164 33
rect 39 30 164 31
rect 39 19 43 30
rect 119 29 164 30
rect 38 18 43 19
rect 38 16 39 18
rect 41 16 43 18
rect 38 15 43 16
rect 38 13 42 15
rect 172 5 177 143
rect 172 3 174 5
rect 176 3 177 5
rect 172 1 177 3
rect 187 -2 191 348
rect 384 310 413 311
rect 264 309 414 310
rect 264 307 265 309
rect 267 307 414 309
rect 264 305 414 307
rect 279 304 386 305
rect 410 290 414 305
rect 410 288 411 290
rect 413 288 414 290
rect 410 286 414 288
rect 534 302 538 303
rect 534 300 535 302
rect 537 300 538 302
rect 534 289 538 300
rect 1020 289 1091 292
rect 534 288 729 289
rect 534 286 726 288
rect 728 286 729 288
rect 534 285 729 286
rect 1020 287 1088 289
rect 1090 287 1091 289
rect 1020 286 1091 287
rect 324 167 335 168
rect 324 166 329 167
rect 324 164 325 166
rect 327 165 329 166
rect 331 165 335 167
rect 327 164 335 165
rect 324 162 335 164
rect 593 89 612 90
rect 593 87 598 89
rect 600 87 603 89
rect 605 87 612 89
rect 593 85 612 87
rect 1020 75 1025 286
rect 548 73 675 75
rect 548 72 672 73
rect 548 70 550 72
rect 552 71 672 72
rect 674 71 675 73
rect 552 70 675 71
rect 548 67 675 70
rect 1019 68 1025 75
rect 269 63 274 64
rect 269 61 270 63
rect 272 61 274 63
rect 269 33 274 61
rect 868 46 879 47
rect 868 44 870 46
rect 872 44 876 46
rect 878 44 879 46
rect 868 43 879 44
rect 196 32 629 33
rect 196 30 197 32
rect 199 30 629 32
rect 196 28 629 30
rect 187 -4 188 -2
rect 190 -4 191 -2
rect 187 -6 191 -4
rect 210 4 214 6
rect 210 2 211 4
rect 213 2 214 4
rect -24 -17 -23 -15
rect -21 -17 -20 -15
rect -24 -18 -20 -17
rect 24 -12 28 -10
rect 24 -14 25 -12
rect 27 -14 28 -12
rect 24 -17 28 -14
rect 24 -19 25 -17
rect 27 -19 28 -17
rect 24 -20 28 -19
rect 210 -43 214 2
rect 235 2 241 4
rect 235 0 237 2
rect 239 0 241 2
rect 235 -1 241 0
rect 210 -45 211 -43
rect 213 -45 214 -43
rect 210 -47 214 -45
rect 237 -46 241 -1
rect 237 -48 238 -46
rect 240 -48 241 -46
rect 252 3 256 4
rect 252 1 253 3
rect 255 1 256 3
rect 252 -45 256 1
rect 269 -39 274 28
rect 625 -7 629 28
rect 1019 5 1024 68
rect 840 3 1024 5
rect 840 1 842 3
rect 844 1 1024 3
rect 840 -1 1024 1
rect 338 -10 520 -8
rect 338 -12 517 -10
rect 519 -12 520 -10
rect 338 -13 520 -12
rect 625 -9 626 -7
rect 628 -9 629 -7
rect 289 -18 342 -13
rect 289 -38 293 -18
rect 346 -22 374 -20
rect 346 -24 347 -22
rect 349 -24 371 -22
rect 373 -24 374 -22
rect 346 -25 374 -24
rect 625 -25 629 -9
rect 324 -31 461 -29
rect 324 -33 327 -31
rect 329 -33 458 -31
rect 460 -33 461 -31
rect 324 -34 461 -33
rect 269 -41 271 -39
rect 273 -41 274 -39
rect 269 -43 274 -41
rect 285 -39 293 -38
rect 285 -41 289 -39
rect 291 -41 293 -39
rect 285 -43 293 -41
rect 300 -40 304 -39
rect 300 -42 301 -40
rect 303 -42 304 -40
rect 252 -47 253 -45
rect 255 -47 256 -45
rect 252 -48 256 -47
rect 162 -58 166 -48
rect 237 -50 241 -48
rect 283 -52 288 -50
rect 283 -54 285 -52
rect 287 -54 288 -52
rect 283 -58 288 -54
rect 162 -59 288 -58
rect 162 -61 163 -59
rect 165 -61 288 -59
rect 162 -63 288 -61
rect 300 -80 304 -42
rect 334 -41 338 -38
rect 334 -43 335 -41
rect 337 -43 338 -41
rect 334 -62 338 -43
rect 334 -64 335 -62
rect 337 -64 338 -62
rect 334 -65 338 -64
<< alu5 >>
rect 16 273 41 274
rect 16 271 17 273
rect 19 271 38 273
rect 40 271 41 273
rect 16 270 41 271
rect -282 167 335 168
rect -282 165 -281 167
rect -279 166 335 167
rect -279 165 325 166
rect -282 164 325 165
rect 327 164 335 166
rect 320 162 335 164
rect -41 120 -37 124
rect -276 89 612 90
rect -276 87 -274 89
rect -272 87 598 89
rect 600 87 612 89
rect -276 86 612 87
rect -34 85 612 86
rect -276 46 873 47
rect -276 44 -274 46
rect -272 44 870 46
rect 872 44 873 46
rect -276 43 873 44
rect -41 1 28 3
rect -41 -1 -40 1
rect -38 -1 28 1
rect -41 -2 28 -1
rect 24 -12 28 -2
rect 24 -14 25 -12
rect 27 -14 28 -12
rect 24 -15 28 -14
<< ptie >>
rect -282 295 -276 297
rect -282 293 -280 295
rect -278 293 -276 295
rect -282 291 -276 293
rect -7 295 -1 297
rect -7 293 -5 295
rect -3 293 -1 295
rect -7 291 -1 293
rect 36 295 42 297
rect 36 293 38 295
rect 40 293 42 295
rect 36 291 42 293
rect 76 295 82 297
rect 76 293 78 295
rect 80 293 82 295
rect 76 291 82 293
rect 295 295 301 297
rect 295 293 297 295
rect 299 293 301 295
rect 295 291 301 293
rect 343 295 349 297
rect 343 293 345 295
rect 347 293 349 295
rect 343 291 349 293
rect 572 295 578 297
rect 572 293 574 295
rect 576 293 578 295
rect 572 291 578 293
rect 620 295 626 297
rect 620 293 622 295
rect 624 293 626 295
rect 620 291 626 293
rect 848 295 854 297
rect 848 293 850 295
rect 852 293 854 295
rect 848 291 854 293
rect 896 295 902 297
rect 896 293 898 295
rect 900 293 902 295
rect 896 291 902 293
rect 1125 295 1131 297
rect 1125 293 1127 295
rect 1129 293 1131 295
rect 1125 291 1131 293
rect -282 283 -276 285
rect -282 281 -280 283
rect -278 281 -276 283
rect -282 279 -276 281
rect -7 283 -1 285
rect -7 281 -5 283
rect -3 281 -1 283
rect -7 279 -1 281
rect 36 283 42 285
rect 36 281 38 283
rect 40 281 42 283
rect 36 279 42 281
rect 76 283 82 285
rect 76 281 78 283
rect 80 281 82 283
rect 76 279 82 281
rect 295 283 301 285
rect 295 281 297 283
rect 299 281 301 283
rect 295 279 301 281
rect 343 283 349 285
rect 343 281 345 283
rect 347 281 349 283
rect 343 279 349 281
rect 572 283 578 285
rect 572 281 574 283
rect 576 281 578 283
rect 572 279 578 281
rect 620 283 626 285
rect 620 281 622 283
rect 624 281 626 283
rect 620 279 626 281
rect 848 283 854 285
rect 848 281 850 283
rect 852 281 854 283
rect 848 279 854 281
rect 896 283 902 285
rect 896 281 898 283
rect 900 281 902 283
rect 896 279 902 281
rect 1125 283 1131 285
rect 1125 281 1127 283
rect 1129 281 1131 283
rect 1125 279 1131 281
rect -282 151 -276 153
rect -282 149 -280 151
rect -278 149 -276 151
rect -282 147 -276 149
rect -7 151 -1 153
rect -7 149 -5 151
rect -3 149 -1 151
rect -7 147 -1 149
rect 36 151 42 153
rect 36 149 38 151
rect 40 149 42 151
rect 36 147 42 149
rect 76 151 82 153
rect 76 149 78 151
rect 80 149 82 151
rect 76 147 82 149
rect 295 151 301 153
rect 295 149 297 151
rect 299 149 301 151
rect 295 147 301 149
rect 343 151 349 153
rect 343 149 345 151
rect 347 149 349 151
rect 343 147 349 149
rect 572 151 578 153
rect 572 149 574 151
rect 576 149 578 151
rect 572 147 578 149
rect 620 151 626 153
rect 620 149 622 151
rect 624 149 626 151
rect 620 147 626 149
rect 848 151 854 153
rect 848 149 850 151
rect 852 149 854 151
rect 848 147 854 149
rect 896 151 902 153
rect 896 149 898 151
rect 900 149 902 151
rect 896 147 902 149
rect 1125 151 1131 153
rect 1125 149 1127 151
rect 1129 149 1131 151
rect 1125 147 1131 149
rect -282 139 -276 141
rect -282 137 -280 139
rect -278 137 -276 139
rect -282 135 -276 137
rect -7 139 -1 141
rect -7 137 -5 139
rect -3 137 -1 139
rect -7 135 -1 137
rect 36 139 42 141
rect 36 137 38 139
rect 40 137 42 139
rect 36 135 42 137
rect 76 139 82 141
rect 76 137 78 139
rect 80 137 82 139
rect 76 135 82 137
rect 295 139 301 141
rect 295 137 297 139
rect 299 137 301 139
rect 295 135 301 137
rect 343 139 349 141
rect 343 137 345 139
rect 347 137 349 139
rect 343 135 349 137
rect 572 139 578 141
rect 572 137 574 139
rect 576 137 578 139
rect 572 135 578 137
rect 620 139 626 141
rect 620 137 622 139
rect 624 137 626 139
rect 620 135 626 137
rect 848 139 854 141
rect 848 137 850 139
rect 852 137 854 139
rect 848 135 854 137
rect 896 139 902 141
rect 896 137 898 139
rect 900 137 902 139
rect 896 135 902 137
rect 1125 139 1131 141
rect 1125 137 1127 139
rect 1129 137 1131 139
rect 1125 135 1131 137
rect -282 7 -276 9
rect -282 5 -280 7
rect -278 5 -276 7
rect -282 3 -276 5
rect -7 7 -1 9
rect -7 5 -5 7
rect -3 5 -1 7
rect -7 3 -1 5
rect 36 7 42 9
rect 36 5 38 7
rect 40 5 42 7
rect 36 3 42 5
rect 76 7 82 9
rect 76 5 78 7
rect 80 5 82 7
rect 76 3 82 5
rect 295 7 301 9
rect 295 5 297 7
rect 299 5 301 7
rect 295 3 301 5
rect 343 7 349 9
rect 343 5 345 7
rect 347 5 349 7
rect 343 3 349 5
rect 572 7 578 9
rect 572 5 574 7
rect 576 5 578 7
rect 572 3 578 5
rect 620 7 626 9
rect 620 5 622 7
rect 624 5 626 7
rect 620 3 626 5
rect 848 7 854 9
rect 848 5 850 7
rect 852 5 854 7
rect 848 3 854 5
rect 896 7 902 9
rect 896 5 898 7
rect 900 5 902 7
rect 896 3 902 5
rect 1125 7 1131 9
rect 1125 5 1127 7
rect 1129 5 1131 7
rect 1125 3 1131 5
rect -155 -4 -149 -2
rect -155 -6 -153 -4
rect -151 -6 -149 -4
rect -155 -8 -149 -6
rect -123 -4 -109 -2
rect -123 -6 -121 -4
rect -119 -6 -113 -4
rect -111 -6 -109 -4
rect -123 -8 -109 -6
rect -103 -4 -97 -2
rect -103 -6 -101 -4
rect -99 -6 -97 -4
rect -103 -8 -97 -6
rect -71 -4 -57 -2
rect -71 -6 -69 -4
rect -67 -6 -61 -4
rect -59 -6 -57 -4
rect -71 -8 -57 -6
rect -51 -4 -45 -2
rect -51 -6 -49 -4
rect -47 -6 -45 -4
rect -51 -8 -45 -6
rect -19 -4 -5 -2
rect -19 -6 -17 -4
rect -15 -6 -9 -4
rect -7 -6 -5 -4
rect -19 -8 -5 -6
rect 1 -4 7 -2
rect 1 -6 3 -4
rect 5 -6 7 -4
rect 1 -8 7 -6
rect 33 -4 47 -2
rect 33 -6 35 -4
rect 37 -6 43 -4
rect 45 -6 47 -4
rect 33 -8 47 -6
rect 53 -4 59 -2
rect 53 -6 55 -4
rect 57 -6 59 -4
rect 53 -8 59 -6
rect 85 -4 99 -2
rect 85 -6 87 -4
rect 89 -6 95 -4
rect 97 -6 99 -4
rect 85 -8 99 -6
rect 106 -4 112 -2
rect 106 -6 108 -4
rect 110 -6 112 -4
rect 106 -8 112 -6
rect 138 -4 152 -2
rect 138 -6 140 -4
rect 142 -6 148 -4
rect 150 -6 152 -4
rect 138 -8 152 -6
rect 163 -4 177 -2
rect 163 -6 165 -4
rect 167 -6 173 -4
rect 175 -6 177 -4
rect 163 -11 177 -6
rect 183 -4 197 -2
rect 183 -6 185 -4
rect 187 -6 193 -4
rect 195 -6 197 -4
rect 183 -11 197 -6
rect 203 -4 217 -2
rect 203 -6 205 -4
rect 207 -6 213 -4
rect 215 -6 217 -4
rect 203 -11 217 -6
rect 225 -4 239 -2
rect 225 -6 227 -4
rect 229 -6 235 -4
rect 237 -6 239 -4
rect 225 -11 239 -6
rect 247 -4 261 -2
rect 247 -6 249 -4
rect 251 -6 257 -4
rect 259 -6 261 -4
rect 247 -11 261 -6
rect 269 -4 283 -2
rect 269 -6 271 -4
rect 273 -6 279 -4
rect 281 -6 283 -4
rect 269 -11 283 -6
rect 294 -4 300 -2
rect 294 -6 296 -4
rect 298 -6 300 -4
rect 294 -8 300 -6
rect 326 -4 340 -2
rect 326 -6 328 -4
rect 330 -6 336 -4
rect 338 -6 340 -4
rect 326 -8 340 -6
rect 347 -4 353 -2
rect 347 -6 349 -4
rect 351 -6 353 -4
rect 347 -8 353 -6
rect 379 -4 393 -2
rect 379 -6 381 -4
rect 383 -6 389 -4
rect 391 -6 393 -4
rect 379 -8 393 -6
rect 399 -4 405 -2
rect 399 -6 401 -4
rect 403 -6 405 -4
rect 399 -8 405 -6
rect 431 -4 445 -2
rect 431 -6 433 -4
rect 435 -6 441 -4
rect 443 -6 445 -4
rect 431 -8 445 -6
rect 451 -4 457 -2
rect 451 -6 453 -4
rect 455 -6 457 -4
rect 451 -8 457 -6
rect 483 -4 497 -2
rect 483 -6 485 -4
rect 487 -6 493 -4
rect 495 -6 497 -4
rect 483 -8 497 -6
rect 503 -4 509 -2
rect 503 -6 505 -4
rect 507 -6 509 -4
rect 503 -8 509 -6
rect 535 -4 549 -2
rect 535 -6 537 -4
rect 539 -6 545 -4
rect 547 -6 549 -4
rect 535 -8 549 -6
rect 558 -4 572 -2
rect 558 -6 560 -4
rect 562 -6 568 -4
rect 570 -6 572 -4
rect 558 -11 572 -6
rect 579 -4 593 -2
rect 579 -6 581 -4
rect 583 -6 589 -4
rect 591 -6 593 -4
rect 579 -11 593 -6
rect 602 -4 608 -2
rect 602 -6 604 -4
rect 606 -6 608 -4
rect 602 -8 608 -6
rect 634 -4 648 -2
rect 634 -6 636 -4
rect 638 -6 644 -4
rect 646 -6 648 -4
rect 634 -8 648 -6
rect 655 -4 661 -2
rect 655 -6 657 -4
rect 659 -6 661 -4
rect 655 -8 661 -6
rect 687 -4 701 -2
rect 687 -6 689 -4
rect 691 -6 697 -4
rect 699 -6 701 -4
rect 687 -8 701 -6
rect 707 -4 713 -2
rect 707 -6 709 -4
rect 711 -6 713 -4
rect 707 -8 713 -6
rect 739 -4 753 -2
rect 739 -6 741 -4
rect 743 -6 749 -4
rect 751 -6 753 -4
rect 739 -8 753 -6
rect 759 -4 765 -2
rect 759 -6 761 -4
rect 763 -6 765 -4
rect 759 -8 765 -6
rect 791 -4 805 -2
rect 791 -6 793 -4
rect 795 -6 801 -4
rect 803 -6 805 -4
rect 791 -8 805 -6
rect 811 -4 817 -2
rect 811 -6 813 -4
rect 815 -6 817 -4
rect 811 -8 817 -6
rect 843 -4 857 -2
rect 843 -6 845 -4
rect 847 -6 853 -4
rect 855 -6 857 -4
rect 843 -8 857 -6
rect 863 -4 869 -2
rect 863 -6 865 -4
rect 867 -6 869 -4
rect 863 -8 869 -6
rect 895 -4 909 -2
rect 895 -6 897 -4
rect 899 -6 905 -4
rect 907 -6 909 -4
rect 895 -8 909 -6
rect 916 -4 922 -2
rect 916 -6 918 -4
rect 920 -6 922 -4
rect 916 -8 922 -6
rect 948 -4 962 -2
rect 948 -6 950 -4
rect 952 -6 958 -4
rect 960 -6 962 -4
rect 948 -8 962 -6
rect 970 -4 976 -2
rect 970 -6 972 -4
rect 974 -6 976 -4
rect 970 -8 976 -6
rect 1002 -4 1016 -2
rect 1002 -6 1004 -4
rect 1006 -6 1012 -4
rect 1014 -6 1016 -4
rect 1002 -8 1016 -6
rect 1025 -4 1031 -2
rect 1025 -6 1027 -4
rect 1029 -6 1031 -4
rect 1025 -8 1031 -6
rect 1057 -4 1071 -2
rect 1057 -6 1059 -4
rect 1061 -6 1067 -4
rect 1069 -6 1071 -4
rect 1057 -8 1071 -6
rect 1078 -4 1084 -2
rect 1078 -6 1080 -4
rect 1082 -6 1084 -4
rect 1078 -8 1084 -6
rect 1110 -4 1124 -2
rect 1110 -6 1112 -4
rect 1114 -6 1120 -4
rect 1122 -6 1124 -4
rect 1110 -8 1124 -6
<< ntie >>
rect -249 355 -243 357
rect -249 353 -247 355
rect -245 353 -243 355
rect -249 351 -243 353
rect -7 355 -1 357
rect -7 353 -5 355
rect -3 353 -1 355
rect -7 351 -1 353
rect 36 355 42 357
rect 36 353 38 355
rect 40 353 42 355
rect 36 351 42 353
rect 76 355 82 357
rect 76 353 78 355
rect 80 353 82 355
rect 76 351 82 353
rect 295 355 301 357
rect 295 353 297 355
rect 299 353 301 355
rect 295 351 301 353
rect 343 355 349 357
rect 343 353 345 355
rect 347 353 349 355
rect 343 351 349 353
rect 572 355 578 357
rect 572 353 574 355
rect 576 353 578 355
rect 572 351 578 353
rect 620 355 626 357
rect 620 353 622 355
rect 624 353 626 355
rect 620 351 626 353
rect 848 355 854 357
rect 848 353 850 355
rect 852 353 854 355
rect 848 351 854 353
rect 896 355 902 357
rect 896 353 898 355
rect 900 353 902 355
rect 896 351 902 353
rect 1125 355 1131 357
rect 1125 353 1127 355
rect 1129 353 1131 355
rect 1125 351 1131 353
rect -249 223 -243 225
rect -249 221 -247 223
rect -245 221 -243 223
rect -249 219 -243 221
rect -7 223 -1 225
rect -7 221 -5 223
rect -3 221 -1 223
rect -7 219 -1 221
rect 36 223 42 225
rect 36 221 38 223
rect 40 221 42 223
rect 36 219 42 221
rect 76 223 82 225
rect 76 221 78 223
rect 80 221 82 223
rect 76 219 82 221
rect 295 223 301 225
rect 295 221 297 223
rect 299 221 301 223
rect 295 219 301 221
rect 343 223 349 225
rect 343 221 345 223
rect 347 221 349 223
rect 343 219 349 221
rect 572 223 578 225
rect 572 221 574 223
rect 576 221 578 223
rect 572 219 578 221
rect 620 223 626 225
rect 620 221 622 223
rect 624 221 626 223
rect 620 219 626 221
rect 848 223 854 225
rect 848 221 850 223
rect 852 221 854 223
rect 848 219 854 221
rect 896 223 902 225
rect 896 221 898 223
rect 900 221 902 223
rect 896 219 902 221
rect 1125 223 1131 225
rect 1125 221 1127 223
rect 1129 221 1131 223
rect 1125 219 1131 221
rect -249 211 -243 213
rect -249 209 -247 211
rect -245 209 -243 211
rect -249 207 -243 209
rect -7 211 -1 213
rect -7 209 -5 211
rect -3 209 -1 211
rect -7 207 -1 209
rect 36 211 42 213
rect 36 209 38 211
rect 40 209 42 211
rect 36 207 42 209
rect 76 211 82 213
rect 76 209 78 211
rect 80 209 82 211
rect 76 207 82 209
rect 295 211 301 213
rect 295 209 297 211
rect 299 209 301 211
rect 295 207 301 209
rect 343 211 349 213
rect 343 209 345 211
rect 347 209 349 211
rect 343 207 349 209
rect 572 211 578 213
rect 572 209 574 211
rect 576 209 578 211
rect 572 207 578 209
rect 620 211 626 213
rect 620 209 622 211
rect 624 209 626 211
rect 620 207 626 209
rect 848 211 854 213
rect 848 209 850 211
rect 852 209 854 211
rect 848 207 854 209
rect 896 211 902 213
rect 896 209 898 211
rect 900 209 902 211
rect 896 207 902 209
rect 1125 211 1131 213
rect 1125 209 1127 211
rect 1129 209 1131 211
rect 1125 207 1131 209
rect -249 79 -243 81
rect -249 77 -247 79
rect -245 77 -243 79
rect -249 75 -243 77
rect -7 79 -1 81
rect -7 77 -5 79
rect -3 77 -1 79
rect -7 75 -1 77
rect 36 79 42 81
rect 36 77 38 79
rect 40 77 42 79
rect 36 75 42 77
rect 76 79 82 81
rect 76 77 78 79
rect 80 77 82 79
rect 76 75 82 77
rect 295 79 301 81
rect 295 77 297 79
rect 299 77 301 79
rect 295 75 301 77
rect 343 79 349 81
rect 343 77 345 79
rect 347 77 349 79
rect 343 75 349 77
rect 572 79 578 81
rect 572 77 574 79
rect 576 77 578 79
rect 572 75 578 77
rect 620 79 626 81
rect 620 77 622 79
rect 624 77 626 79
rect 620 75 626 77
rect 848 79 854 81
rect 848 77 850 79
rect 852 77 854 79
rect 848 75 854 77
rect 896 79 902 81
rect 896 77 898 79
rect 900 77 902 79
rect 896 75 902 77
rect 1125 79 1131 81
rect 1125 77 1127 79
rect 1129 77 1131 79
rect 1125 75 1131 77
rect -249 67 -243 69
rect -249 65 -247 67
rect -245 65 -243 67
rect -249 63 -243 65
rect -7 67 -1 69
rect -7 65 -5 67
rect -3 65 -1 67
rect -7 63 -1 65
rect 36 67 42 69
rect 36 65 38 67
rect 40 65 42 67
rect 36 63 42 65
rect 76 67 82 69
rect 76 65 78 67
rect 80 65 82 67
rect 76 63 82 65
rect 295 67 301 69
rect 295 65 297 67
rect 299 65 301 67
rect 295 63 301 65
rect 343 67 349 69
rect 343 65 345 67
rect 347 65 349 67
rect 343 63 349 65
rect 572 67 578 69
rect 572 65 574 67
rect 576 65 578 67
rect 572 63 578 65
rect 620 67 626 69
rect 620 65 622 67
rect 624 65 626 67
rect 620 63 626 65
rect 848 67 854 69
rect 848 65 850 67
rect 852 65 854 67
rect 848 63 854 65
rect 896 67 902 69
rect 896 65 898 67
rect 900 65 902 67
rect 896 63 902 65
rect 1125 67 1131 69
rect 1125 65 1127 67
rect 1129 65 1131 67
rect 1125 63 1131 65
rect -135 -64 -129 -62
rect -135 -66 -133 -64
rect -131 -66 -129 -64
rect -135 -68 -129 -66
rect -83 -64 -77 -62
rect -83 -66 -81 -64
rect -79 -66 -77 -64
rect -83 -68 -77 -66
rect -31 -64 -25 -62
rect -31 -66 -29 -64
rect -27 -66 -25 -64
rect -31 -68 -25 -66
rect 21 -64 27 -62
rect 21 -66 23 -64
rect 25 -66 27 -64
rect 21 -68 27 -66
rect 73 -64 79 -62
rect 73 -66 75 -64
rect 77 -66 79 -64
rect 73 -68 79 -66
rect 126 -64 132 -62
rect 126 -66 128 -64
rect 130 -66 132 -64
rect 126 -68 132 -66
rect 172 -64 178 -61
rect 172 -66 174 -64
rect 176 -66 178 -64
rect 172 -68 178 -66
rect 192 -64 198 -61
rect 192 -66 194 -64
rect 196 -66 198 -64
rect 192 -68 198 -66
rect 212 -64 218 -61
rect 212 -66 214 -64
rect 216 -66 218 -64
rect 212 -68 218 -66
rect 234 -64 240 -61
rect 234 -66 236 -64
rect 238 -66 240 -64
rect 234 -68 240 -66
rect 256 -64 262 -61
rect 256 -66 258 -64
rect 260 -66 262 -64
rect 256 -68 262 -66
rect 278 -64 284 -61
rect 278 -66 280 -64
rect 282 -66 284 -64
rect 278 -68 284 -66
rect 314 -64 320 -62
rect 314 -66 316 -64
rect 318 -66 320 -64
rect 314 -68 320 -66
rect 367 -64 373 -62
rect 367 -66 369 -64
rect 371 -66 373 -64
rect 367 -68 373 -66
rect 419 -64 425 -62
rect 419 -66 421 -64
rect 423 -66 425 -64
rect 419 -68 425 -66
rect 471 -64 477 -62
rect 471 -66 473 -64
rect 475 -66 477 -64
rect 471 -68 477 -66
rect 523 -64 529 -62
rect 523 -66 525 -64
rect 527 -66 529 -64
rect 523 -68 529 -66
rect 567 -64 573 -61
rect 567 -66 569 -64
rect 571 -66 573 -64
rect 567 -68 573 -66
rect 588 -64 594 -61
rect 588 -66 590 -64
rect 592 -66 594 -64
rect 588 -68 594 -66
rect 622 -64 628 -62
rect 622 -66 624 -64
rect 626 -66 628 -64
rect 622 -68 628 -66
rect 675 -64 681 -62
rect 675 -66 677 -64
rect 679 -66 681 -64
rect 675 -68 681 -66
rect 727 -64 733 -62
rect 727 -66 729 -64
rect 731 -66 733 -64
rect 727 -68 733 -66
rect 779 -64 785 -62
rect 779 -66 781 -64
rect 783 -66 785 -64
rect 779 -68 785 -66
rect 831 -64 837 -62
rect 831 -66 833 -64
rect 835 -66 837 -64
rect 831 -68 837 -66
rect 883 -64 889 -62
rect 883 -66 885 -64
rect 887 -66 889 -64
rect 883 -68 889 -66
rect 936 -64 942 -62
rect 936 -66 938 -64
rect 940 -66 942 -64
rect 936 -68 942 -66
rect 990 -64 996 -62
rect 990 -66 992 -64
rect 994 -66 996 -64
rect 990 -68 996 -66
rect 1045 -64 1051 -62
rect 1045 -66 1047 -64
rect 1049 -66 1051 -64
rect 1045 -68 1051 -66
rect 1098 -64 1104 -62
rect 1098 -66 1100 -64
rect 1102 -66 1104 -64
rect 1098 -68 1104 -66
<< nmos >>
rect -276 305 -274 314
rect -260 300 -258 309
rect -250 300 -248 309
rect -240 297 -238 309
rect -233 297 -231 309
rect -208 294 -206 307
rect -198 297 -196 307
rect -188 300 -186 314
rect -178 300 -176 314
rect -158 294 -156 314
rect -151 294 -149 314
rect -140 294 -138 308
rect -118 294 -116 308
rect -107 294 -105 314
rect -100 294 -98 314
rect -80 300 -78 314
rect -70 300 -68 314
rect -29 308 -27 314
rect -19 308 -17 314
rect -60 297 -58 307
rect -50 294 -48 307
rect -9 305 -7 314
rect 14 301 16 312
rect 21 301 23 312
rect 34 303 36 312
rect 54 301 56 312
rect 61 301 63 312
rect 74 303 76 312
rect 94 294 96 307
rect 104 297 106 307
rect 114 300 116 314
rect 124 300 126 314
rect 144 294 146 314
rect 151 294 153 314
rect 162 294 164 308
rect 184 294 186 308
rect 195 294 197 314
rect 202 294 204 314
rect 222 300 224 314
rect 232 300 234 314
rect 273 308 275 314
rect 283 308 285 314
rect 242 297 244 307
rect 252 294 254 307
rect 293 305 295 314
rect 321 301 323 312
rect 328 301 330 312
rect 341 303 343 312
rect 371 294 373 307
rect 381 297 383 307
rect 391 300 393 314
rect 401 300 403 314
rect 421 294 423 314
rect 428 294 430 314
rect 439 294 441 308
rect 461 294 463 308
rect 472 294 474 314
rect 479 294 481 314
rect 499 300 501 314
rect 509 300 511 314
rect 550 308 552 314
rect 560 308 562 314
rect 519 297 521 307
rect 529 294 531 307
rect 570 305 572 314
rect 598 301 600 312
rect 605 301 607 312
rect 618 303 620 312
rect 647 294 649 307
rect 657 297 659 307
rect 667 300 669 314
rect 677 300 679 314
rect 697 294 699 314
rect 704 294 706 314
rect 715 294 717 308
rect 737 294 739 308
rect 748 294 750 314
rect 755 294 757 314
rect 775 300 777 314
rect 785 300 787 314
rect 826 308 828 314
rect 836 308 838 314
rect 795 297 797 307
rect 805 294 807 307
rect 846 305 848 314
rect 874 301 876 312
rect 881 301 883 312
rect 894 303 896 312
rect 924 294 926 307
rect 934 297 936 307
rect 944 300 946 314
rect 954 300 956 314
rect 974 294 976 314
rect 981 294 983 314
rect 992 294 994 308
rect 1014 294 1016 308
rect 1025 294 1027 314
rect 1032 294 1034 314
rect 1052 300 1054 314
rect 1062 300 1064 314
rect 1103 308 1105 314
rect 1113 308 1115 314
rect 1072 297 1074 307
rect 1082 294 1084 307
rect 1123 305 1125 314
rect -276 262 -274 271
rect -260 267 -258 276
rect -250 267 -248 276
rect -240 267 -238 279
rect -233 267 -231 279
rect -208 269 -206 282
rect -198 269 -196 279
rect -188 262 -186 276
rect -178 262 -176 276
rect -158 262 -156 282
rect -151 262 -149 282
rect -140 268 -138 282
rect -118 268 -116 282
rect -107 262 -105 282
rect -100 262 -98 282
rect -80 262 -78 276
rect -70 262 -68 276
rect -60 269 -58 279
rect -50 269 -48 282
rect -29 262 -27 268
rect -19 262 -17 268
rect -9 262 -7 271
rect 14 264 16 275
rect 21 264 23 275
rect 34 264 36 273
rect 54 264 56 275
rect 61 264 63 275
rect 74 264 76 273
rect 94 269 96 282
rect 104 269 106 279
rect 114 262 116 276
rect 124 262 126 276
rect 144 262 146 282
rect 151 262 153 282
rect 162 268 164 282
rect 184 268 186 282
rect 195 262 197 282
rect 202 262 204 282
rect 222 262 224 276
rect 232 262 234 276
rect 242 269 244 279
rect 252 269 254 282
rect 273 262 275 268
rect 283 262 285 268
rect 293 262 295 271
rect 321 264 323 275
rect 328 264 330 275
rect 341 264 343 273
rect 371 269 373 282
rect 381 269 383 279
rect 391 262 393 276
rect 401 262 403 276
rect 421 262 423 282
rect 428 262 430 282
rect 439 268 441 282
rect 461 268 463 282
rect 472 262 474 282
rect 479 262 481 282
rect 499 262 501 276
rect 509 262 511 276
rect 519 269 521 279
rect 529 269 531 282
rect 550 262 552 268
rect 560 262 562 268
rect 570 262 572 271
rect 598 264 600 275
rect 605 264 607 275
rect 618 264 620 273
rect 647 269 649 282
rect 657 269 659 279
rect 667 262 669 276
rect 677 262 679 276
rect 697 262 699 282
rect 704 262 706 282
rect 715 268 717 282
rect 737 268 739 282
rect 748 262 750 282
rect 755 262 757 282
rect 775 262 777 276
rect 785 262 787 276
rect 795 269 797 279
rect 805 269 807 282
rect 826 262 828 268
rect 836 262 838 268
rect 846 262 848 271
rect 874 264 876 275
rect 881 264 883 275
rect 894 264 896 273
rect 924 269 926 282
rect 934 269 936 279
rect 944 262 946 276
rect 954 262 956 276
rect 974 262 976 282
rect 981 262 983 282
rect 992 268 994 282
rect 1014 268 1016 282
rect 1025 262 1027 282
rect 1032 262 1034 282
rect 1052 262 1054 276
rect 1062 262 1064 276
rect 1072 269 1074 279
rect 1082 269 1084 282
rect 1103 262 1105 268
rect 1113 262 1115 268
rect 1123 262 1125 271
rect -276 161 -274 170
rect -260 156 -258 165
rect -250 156 -248 165
rect -240 153 -238 165
rect -233 153 -231 165
rect -208 150 -206 163
rect -198 153 -196 163
rect -188 156 -186 170
rect -178 156 -176 170
rect -158 150 -156 170
rect -151 150 -149 170
rect -140 150 -138 164
rect -118 150 -116 164
rect -107 150 -105 170
rect -100 150 -98 170
rect -80 156 -78 170
rect -70 156 -68 170
rect -29 164 -27 170
rect -19 164 -17 170
rect -60 153 -58 163
rect -50 150 -48 163
rect -9 161 -7 170
rect 14 157 16 168
rect 21 157 23 168
rect 34 159 36 168
rect 54 157 56 168
rect 61 157 63 168
rect 74 159 76 168
rect 94 150 96 163
rect 104 153 106 163
rect 114 156 116 170
rect 124 156 126 170
rect 144 150 146 170
rect 151 150 153 170
rect 162 150 164 164
rect 184 150 186 164
rect 195 150 197 170
rect 202 150 204 170
rect 222 156 224 170
rect 232 156 234 170
rect 273 164 275 170
rect 283 164 285 170
rect 242 153 244 163
rect 252 150 254 163
rect 293 161 295 170
rect 321 157 323 168
rect 328 157 330 168
rect 341 159 343 168
rect 371 150 373 163
rect 381 153 383 163
rect 391 156 393 170
rect 401 156 403 170
rect 421 150 423 170
rect 428 150 430 170
rect 439 150 441 164
rect 461 150 463 164
rect 472 150 474 170
rect 479 150 481 170
rect 499 156 501 170
rect 509 156 511 170
rect 550 164 552 170
rect 560 164 562 170
rect 519 153 521 163
rect 529 150 531 163
rect 570 161 572 170
rect 598 157 600 168
rect 605 157 607 168
rect 618 159 620 168
rect 647 150 649 163
rect 657 153 659 163
rect 667 156 669 170
rect 677 156 679 170
rect 697 150 699 170
rect 704 150 706 170
rect 715 150 717 164
rect 737 150 739 164
rect 748 150 750 170
rect 755 150 757 170
rect 775 156 777 170
rect 785 156 787 170
rect 826 164 828 170
rect 836 164 838 170
rect 795 153 797 163
rect 805 150 807 163
rect 846 161 848 170
rect 874 157 876 168
rect 881 157 883 168
rect 894 159 896 168
rect 924 150 926 163
rect 934 153 936 163
rect 944 156 946 170
rect 954 156 956 170
rect 974 150 976 170
rect 981 150 983 170
rect 992 150 994 164
rect 1014 150 1016 164
rect 1025 150 1027 170
rect 1032 150 1034 170
rect 1052 156 1054 170
rect 1062 156 1064 170
rect 1103 164 1105 170
rect 1113 164 1115 170
rect 1072 153 1074 163
rect 1082 150 1084 163
rect 1123 161 1125 170
rect -276 118 -274 127
rect -260 123 -258 132
rect -250 123 -248 132
rect -240 123 -238 135
rect -233 123 -231 135
rect -208 125 -206 138
rect -198 125 -196 135
rect -188 118 -186 132
rect -178 118 -176 132
rect -158 118 -156 138
rect -151 118 -149 138
rect -140 124 -138 138
rect -118 124 -116 138
rect -107 118 -105 138
rect -100 118 -98 138
rect -80 118 -78 132
rect -70 118 -68 132
rect -60 125 -58 135
rect -50 125 -48 138
rect -29 118 -27 124
rect -19 118 -17 124
rect -9 118 -7 127
rect 14 120 16 131
rect 21 120 23 131
rect 34 120 36 129
rect 54 120 56 131
rect 61 120 63 131
rect 74 120 76 129
rect 94 125 96 138
rect 104 125 106 135
rect 114 118 116 132
rect 124 118 126 132
rect 144 118 146 138
rect 151 118 153 138
rect 162 124 164 138
rect 184 124 186 138
rect 195 118 197 138
rect 202 118 204 138
rect 222 118 224 132
rect 232 118 234 132
rect 242 125 244 135
rect 252 125 254 138
rect 273 118 275 124
rect 283 118 285 124
rect 293 118 295 127
rect 321 120 323 131
rect 328 120 330 131
rect 341 120 343 129
rect 371 125 373 138
rect 381 125 383 135
rect 391 118 393 132
rect 401 118 403 132
rect 421 118 423 138
rect 428 118 430 138
rect 439 124 441 138
rect 461 124 463 138
rect 472 118 474 138
rect 479 118 481 138
rect 499 118 501 132
rect 509 118 511 132
rect 519 125 521 135
rect 529 125 531 138
rect 550 118 552 124
rect 560 118 562 124
rect 570 118 572 127
rect 598 120 600 131
rect 605 120 607 131
rect 618 120 620 129
rect 647 125 649 138
rect 657 125 659 135
rect 667 118 669 132
rect 677 118 679 132
rect 697 118 699 138
rect 704 118 706 138
rect 715 124 717 138
rect 737 124 739 138
rect 748 118 750 138
rect 755 118 757 138
rect 775 118 777 132
rect 785 118 787 132
rect 795 125 797 135
rect 805 125 807 138
rect 826 118 828 124
rect 836 118 838 124
rect 846 118 848 127
rect 874 120 876 131
rect 881 120 883 131
rect 894 120 896 129
rect 924 125 926 138
rect 934 125 936 135
rect 944 118 946 132
rect 954 118 956 132
rect 974 118 976 138
rect 981 118 983 138
rect 992 124 994 138
rect 1014 124 1016 138
rect 1025 118 1027 138
rect 1032 118 1034 138
rect 1052 118 1054 132
rect 1062 118 1064 132
rect 1072 125 1074 135
rect 1082 125 1084 138
rect 1103 118 1105 124
rect 1113 118 1115 124
rect 1123 118 1125 127
rect -276 17 -274 26
rect -260 12 -258 21
rect -250 12 -248 21
rect -240 9 -238 21
rect -233 9 -231 21
rect -208 6 -206 19
rect -198 9 -196 19
rect -188 12 -186 26
rect -178 12 -176 26
rect -158 6 -156 26
rect -151 6 -149 26
rect -140 6 -138 20
rect -118 6 -116 20
rect -107 6 -105 26
rect -100 6 -98 26
rect -80 12 -78 26
rect -70 12 -68 26
rect -29 20 -27 26
rect -19 20 -17 26
rect -60 9 -58 19
rect -50 6 -48 19
rect -9 17 -7 26
rect 14 13 16 24
rect 21 13 23 24
rect 34 15 36 24
rect 54 13 56 24
rect 61 13 63 24
rect 74 15 76 24
rect 94 6 96 19
rect 104 9 106 19
rect 114 12 116 26
rect 124 12 126 26
rect 144 6 146 26
rect 151 6 153 26
rect 162 6 164 20
rect 184 6 186 20
rect 195 6 197 26
rect 202 6 204 26
rect 222 12 224 26
rect 232 12 234 26
rect 273 20 275 26
rect 283 20 285 26
rect 242 9 244 19
rect 252 6 254 19
rect 293 17 295 26
rect 321 13 323 24
rect 328 13 330 24
rect 341 15 343 24
rect 371 6 373 19
rect 381 9 383 19
rect 391 12 393 26
rect 401 12 403 26
rect 421 6 423 26
rect 428 6 430 26
rect 439 6 441 20
rect 461 6 463 20
rect 472 6 474 26
rect 479 6 481 26
rect 499 12 501 26
rect 509 12 511 26
rect 550 20 552 26
rect 560 20 562 26
rect 519 9 521 19
rect 529 6 531 19
rect 570 17 572 26
rect 598 13 600 24
rect 605 13 607 24
rect 618 15 620 24
rect 647 6 649 19
rect 657 9 659 19
rect 667 12 669 26
rect 677 12 679 26
rect 697 6 699 26
rect 704 6 706 26
rect 715 6 717 20
rect 737 6 739 20
rect 748 6 750 26
rect 755 6 757 26
rect 775 12 777 26
rect 785 12 787 26
rect 826 20 828 26
rect 836 20 838 26
rect 795 9 797 19
rect 805 6 807 19
rect 846 17 848 26
rect 874 13 876 24
rect 881 13 883 24
rect 894 15 896 24
rect 924 6 926 19
rect 934 9 936 19
rect 944 12 946 26
rect 954 12 956 26
rect 974 6 976 26
rect 981 6 983 26
rect 992 6 994 20
rect 1014 6 1016 20
rect 1025 6 1027 26
rect 1032 6 1034 26
rect 1052 12 1054 26
rect 1062 12 1064 26
rect 1103 20 1105 26
rect 1113 20 1115 26
rect 1072 9 1074 19
rect 1082 6 1084 19
rect 1123 17 1125 26
rect -149 -25 -147 -19
rect -134 -25 -132 -14
rect -127 -25 -125 -14
rect -120 -25 -118 -14
rect -97 -25 -95 -19
rect -82 -25 -80 -14
rect -75 -25 -73 -14
rect -68 -25 -66 -14
rect -45 -25 -43 -19
rect -30 -25 -28 -14
rect -23 -25 -21 -14
rect -16 -25 -14 -14
rect 7 -25 9 -19
rect 22 -25 24 -14
rect 29 -25 31 -14
rect 36 -25 38 -14
rect 59 -25 61 -19
rect 74 -25 76 -14
rect 81 -25 83 -14
rect 88 -25 90 -14
rect 112 -25 114 -19
rect 127 -25 129 -14
rect 134 -25 136 -14
rect 141 -25 143 -14
rect 169 -25 171 -19
rect 189 -25 191 -19
rect 209 -25 211 -19
rect 231 -25 233 -19
rect 253 -25 255 -19
rect 275 -25 277 -19
rect 300 -25 302 -19
rect 315 -25 317 -14
rect 322 -25 324 -14
rect 329 -25 331 -14
rect 353 -25 355 -19
rect 368 -25 370 -14
rect 375 -25 377 -14
rect 382 -25 384 -14
rect 405 -25 407 -19
rect 420 -25 422 -14
rect 427 -25 429 -14
rect 434 -25 436 -14
rect 457 -25 459 -19
rect 472 -25 474 -14
rect 479 -25 481 -14
rect 486 -25 488 -14
rect 509 -25 511 -19
rect 524 -25 526 -14
rect 531 -25 533 -14
rect 538 -25 540 -14
rect 564 -25 566 -19
rect 585 -25 587 -19
rect 608 -25 610 -19
rect 623 -25 625 -14
rect 630 -25 632 -14
rect 637 -25 639 -14
rect 661 -25 663 -19
rect 676 -25 678 -14
rect 683 -25 685 -14
rect 690 -25 692 -14
rect 713 -25 715 -19
rect 728 -25 730 -14
rect 735 -25 737 -14
rect 742 -25 744 -14
rect 765 -25 767 -19
rect 780 -25 782 -14
rect 787 -25 789 -14
rect 794 -25 796 -14
rect 817 -25 819 -19
rect 832 -25 834 -14
rect 839 -25 841 -14
rect 846 -25 848 -14
rect 869 -25 871 -19
rect 884 -25 886 -14
rect 891 -25 893 -14
rect 898 -25 900 -14
rect 922 -25 924 -19
rect 937 -25 939 -14
rect 944 -25 946 -14
rect 951 -25 953 -14
rect 976 -25 978 -19
rect 991 -25 993 -14
rect 998 -25 1000 -14
rect 1005 -25 1007 -14
rect 1031 -25 1033 -19
rect 1046 -25 1048 -14
rect 1053 -25 1055 -14
rect 1060 -25 1062 -14
rect 1084 -25 1086 -19
rect 1099 -25 1101 -14
rect 1106 -25 1108 -14
rect 1113 -25 1115 -14
<< pmos >>
rect -268 327 -266 354
rect -252 327 -250 345
rect -242 327 -240 345
rect -232 327 -230 354
rect -208 329 -206 354
rect -195 329 -193 342
rect -185 326 -183 351
rect -178 326 -176 351
rect -160 326 -158 354
rect -150 326 -148 354
rect -140 326 -138 354
rect -118 326 -116 354
rect -108 326 -106 354
rect -98 326 -96 354
rect -80 326 -78 351
rect -73 326 -71 351
rect -63 329 -61 342
rect -50 329 -48 354
rect -29 333 -27 354
rect -22 333 -20 354
rect -9 326 -7 344
rect 14 334 16 347
rect 24 334 26 347
rect 34 327 36 345
rect 54 334 56 347
rect 64 334 66 347
rect 74 327 76 345
rect 94 329 96 354
rect 107 329 109 342
rect 117 326 119 351
rect 124 326 126 351
rect 142 326 144 354
rect 152 326 154 354
rect 162 326 164 354
rect 184 326 186 354
rect 194 326 196 354
rect 204 326 206 354
rect 222 326 224 351
rect 229 326 231 351
rect 239 329 241 342
rect 252 329 254 354
rect 273 333 275 354
rect 280 333 282 354
rect 293 326 295 344
rect 321 334 323 347
rect 331 334 333 347
rect 341 327 343 345
rect 371 329 373 354
rect 384 329 386 342
rect 394 326 396 351
rect 401 326 403 351
rect 419 326 421 354
rect 429 326 431 354
rect 439 326 441 354
rect 461 326 463 354
rect 471 326 473 354
rect 481 326 483 354
rect 499 326 501 351
rect 506 326 508 351
rect 516 329 518 342
rect 529 329 531 354
rect 550 333 552 354
rect 557 333 559 354
rect 570 326 572 344
rect 598 334 600 347
rect 608 334 610 347
rect 618 327 620 345
rect 647 329 649 354
rect 660 329 662 342
rect 670 326 672 351
rect 677 326 679 351
rect 695 326 697 354
rect 705 326 707 354
rect 715 326 717 354
rect 737 326 739 354
rect 747 326 749 354
rect 757 326 759 354
rect 775 326 777 351
rect 782 326 784 351
rect 792 329 794 342
rect 805 329 807 354
rect 826 333 828 354
rect 833 333 835 354
rect 846 326 848 344
rect 874 334 876 347
rect 884 334 886 347
rect 894 327 896 345
rect 924 329 926 354
rect 937 329 939 342
rect 947 326 949 351
rect 954 326 956 351
rect 972 326 974 354
rect 982 326 984 354
rect 992 326 994 354
rect 1014 326 1016 354
rect 1024 326 1026 354
rect 1034 326 1036 354
rect 1052 326 1054 351
rect 1059 326 1061 351
rect 1069 329 1071 342
rect 1082 329 1084 354
rect 1103 333 1105 354
rect 1110 333 1112 354
rect 1123 326 1125 344
rect -268 222 -266 249
rect -252 231 -250 249
rect -242 231 -240 249
rect -232 222 -230 249
rect -208 222 -206 247
rect -195 234 -193 247
rect -185 225 -183 250
rect -178 225 -176 250
rect -160 222 -158 250
rect -150 222 -148 250
rect -140 222 -138 250
rect -118 222 -116 250
rect -108 222 -106 250
rect -98 222 -96 250
rect -80 225 -78 250
rect -73 225 -71 250
rect -63 234 -61 247
rect -50 222 -48 247
rect -29 222 -27 243
rect -22 222 -20 243
rect -9 232 -7 250
rect 14 229 16 242
rect 24 229 26 242
rect 34 231 36 249
rect 54 229 56 242
rect 64 229 66 242
rect 74 231 76 249
rect 94 222 96 247
rect 107 234 109 247
rect 117 225 119 250
rect 124 225 126 250
rect 142 222 144 250
rect 152 222 154 250
rect 162 222 164 250
rect 184 222 186 250
rect 194 222 196 250
rect 204 222 206 250
rect 222 225 224 250
rect 229 225 231 250
rect 239 234 241 247
rect 252 222 254 247
rect 273 222 275 243
rect 280 222 282 243
rect 293 232 295 250
rect 321 229 323 242
rect 331 229 333 242
rect 341 231 343 249
rect 371 222 373 247
rect 384 234 386 247
rect 394 225 396 250
rect 401 225 403 250
rect 419 222 421 250
rect 429 222 431 250
rect 439 222 441 250
rect 461 222 463 250
rect 471 222 473 250
rect 481 222 483 250
rect 499 225 501 250
rect 506 225 508 250
rect 516 234 518 247
rect 529 222 531 247
rect 550 222 552 243
rect 557 222 559 243
rect 570 232 572 250
rect 598 229 600 242
rect 608 229 610 242
rect 618 231 620 249
rect 647 222 649 247
rect 660 234 662 247
rect 670 225 672 250
rect 677 225 679 250
rect 695 222 697 250
rect 705 222 707 250
rect 715 222 717 250
rect 737 222 739 250
rect 747 222 749 250
rect 757 222 759 250
rect 775 225 777 250
rect 782 225 784 250
rect 792 234 794 247
rect 805 222 807 247
rect 826 222 828 243
rect 833 222 835 243
rect 846 232 848 250
rect 874 229 876 242
rect 884 229 886 242
rect 894 231 896 249
rect 924 222 926 247
rect 937 234 939 247
rect 947 225 949 250
rect 954 225 956 250
rect 972 222 974 250
rect 982 222 984 250
rect 992 222 994 250
rect 1014 222 1016 250
rect 1024 222 1026 250
rect 1034 222 1036 250
rect 1052 225 1054 250
rect 1059 225 1061 250
rect 1069 234 1071 247
rect 1082 222 1084 247
rect 1103 222 1105 243
rect 1110 222 1112 243
rect 1123 232 1125 250
rect -268 183 -266 210
rect -252 183 -250 201
rect -242 183 -240 201
rect -232 183 -230 210
rect -208 185 -206 210
rect -195 185 -193 198
rect -185 182 -183 207
rect -178 182 -176 207
rect -160 182 -158 210
rect -150 182 -148 210
rect -140 182 -138 210
rect -118 182 -116 210
rect -108 182 -106 210
rect -98 182 -96 210
rect -80 182 -78 207
rect -73 182 -71 207
rect -63 185 -61 198
rect -50 185 -48 210
rect -29 189 -27 210
rect -22 189 -20 210
rect -9 182 -7 200
rect 14 190 16 203
rect 24 190 26 203
rect 34 183 36 201
rect 54 190 56 203
rect 64 190 66 203
rect 74 183 76 201
rect 94 185 96 210
rect 107 185 109 198
rect 117 182 119 207
rect 124 182 126 207
rect 142 182 144 210
rect 152 182 154 210
rect 162 182 164 210
rect 184 182 186 210
rect 194 182 196 210
rect 204 182 206 210
rect 222 182 224 207
rect 229 182 231 207
rect 239 185 241 198
rect 252 185 254 210
rect 273 189 275 210
rect 280 189 282 210
rect 293 182 295 200
rect 321 190 323 203
rect 331 190 333 203
rect 341 183 343 201
rect 371 185 373 210
rect 384 185 386 198
rect 394 182 396 207
rect 401 182 403 207
rect 419 182 421 210
rect 429 182 431 210
rect 439 182 441 210
rect 461 182 463 210
rect 471 182 473 210
rect 481 182 483 210
rect 499 182 501 207
rect 506 182 508 207
rect 516 185 518 198
rect 529 185 531 210
rect 550 189 552 210
rect 557 189 559 210
rect 570 182 572 200
rect 598 190 600 203
rect 608 190 610 203
rect 618 183 620 201
rect 647 185 649 210
rect 660 185 662 198
rect 670 182 672 207
rect 677 182 679 207
rect 695 182 697 210
rect 705 182 707 210
rect 715 182 717 210
rect 737 182 739 210
rect 747 182 749 210
rect 757 182 759 210
rect 775 182 777 207
rect 782 182 784 207
rect 792 185 794 198
rect 805 185 807 210
rect 826 189 828 210
rect 833 189 835 210
rect 846 182 848 200
rect 874 190 876 203
rect 884 190 886 203
rect 894 183 896 201
rect 924 185 926 210
rect 937 185 939 198
rect 947 182 949 207
rect 954 182 956 207
rect 972 182 974 210
rect 982 182 984 210
rect 992 182 994 210
rect 1014 182 1016 210
rect 1024 182 1026 210
rect 1034 182 1036 210
rect 1052 182 1054 207
rect 1059 182 1061 207
rect 1069 185 1071 198
rect 1082 185 1084 210
rect 1103 189 1105 210
rect 1110 189 1112 210
rect 1123 182 1125 200
rect -268 78 -266 105
rect -252 87 -250 105
rect -242 87 -240 105
rect -232 78 -230 105
rect -208 78 -206 103
rect -195 90 -193 103
rect -185 81 -183 106
rect -178 81 -176 106
rect -160 78 -158 106
rect -150 78 -148 106
rect -140 78 -138 106
rect -118 78 -116 106
rect -108 78 -106 106
rect -98 78 -96 106
rect -80 81 -78 106
rect -73 81 -71 106
rect -63 90 -61 103
rect -50 78 -48 103
rect -29 78 -27 99
rect -22 78 -20 99
rect -9 88 -7 106
rect 14 85 16 98
rect 24 85 26 98
rect 34 87 36 105
rect 54 85 56 98
rect 64 85 66 98
rect 74 87 76 105
rect 94 78 96 103
rect 107 90 109 103
rect 117 81 119 106
rect 124 81 126 106
rect 142 78 144 106
rect 152 78 154 106
rect 162 78 164 106
rect 184 78 186 106
rect 194 78 196 106
rect 204 78 206 106
rect 222 81 224 106
rect 229 81 231 106
rect 239 90 241 103
rect 252 78 254 103
rect 273 78 275 99
rect 280 78 282 99
rect 293 88 295 106
rect 321 85 323 98
rect 331 85 333 98
rect 341 87 343 105
rect 371 78 373 103
rect 384 90 386 103
rect 394 81 396 106
rect 401 81 403 106
rect 419 78 421 106
rect 429 78 431 106
rect 439 78 441 106
rect 461 78 463 106
rect 471 78 473 106
rect 481 78 483 106
rect 499 81 501 106
rect 506 81 508 106
rect 516 90 518 103
rect 529 78 531 103
rect 550 78 552 99
rect 557 78 559 99
rect 570 88 572 106
rect 598 85 600 98
rect 608 85 610 98
rect 618 87 620 105
rect 647 78 649 103
rect 660 90 662 103
rect 670 81 672 106
rect 677 81 679 106
rect 695 78 697 106
rect 705 78 707 106
rect 715 78 717 106
rect 737 78 739 106
rect 747 78 749 106
rect 757 78 759 106
rect 775 81 777 106
rect 782 81 784 106
rect 792 90 794 103
rect 805 78 807 103
rect 826 78 828 99
rect 833 78 835 99
rect 846 88 848 106
rect 874 85 876 98
rect 884 85 886 98
rect 894 87 896 105
rect 924 78 926 103
rect 937 90 939 103
rect 947 81 949 106
rect 954 81 956 106
rect 972 78 974 106
rect 982 78 984 106
rect 992 78 994 106
rect 1014 78 1016 106
rect 1024 78 1026 106
rect 1034 78 1036 106
rect 1052 81 1054 106
rect 1059 81 1061 106
rect 1069 90 1071 103
rect 1082 78 1084 103
rect 1103 78 1105 99
rect 1110 78 1112 99
rect 1123 88 1125 106
rect -268 39 -266 66
rect -252 39 -250 57
rect -242 39 -240 57
rect -232 39 -230 66
rect -208 41 -206 66
rect -195 41 -193 54
rect -185 38 -183 63
rect -178 38 -176 63
rect -160 38 -158 66
rect -150 38 -148 66
rect -140 38 -138 66
rect -118 38 -116 66
rect -108 38 -106 66
rect -98 38 -96 66
rect -80 38 -78 63
rect -73 38 -71 63
rect -63 41 -61 54
rect -50 41 -48 66
rect -29 45 -27 66
rect -22 45 -20 66
rect -9 38 -7 56
rect 14 46 16 59
rect 24 46 26 59
rect 34 39 36 57
rect 54 46 56 59
rect 64 46 66 59
rect 74 39 76 57
rect 94 41 96 66
rect 107 41 109 54
rect 117 38 119 63
rect 124 38 126 63
rect 142 38 144 66
rect 152 38 154 66
rect 162 38 164 66
rect 184 38 186 66
rect 194 38 196 66
rect 204 38 206 66
rect 222 38 224 63
rect 229 38 231 63
rect 239 41 241 54
rect 252 41 254 66
rect 273 45 275 66
rect 280 45 282 66
rect 293 38 295 56
rect 321 46 323 59
rect 331 46 333 59
rect 341 39 343 57
rect 371 41 373 66
rect 384 41 386 54
rect 394 38 396 63
rect 401 38 403 63
rect 419 38 421 66
rect 429 38 431 66
rect 439 38 441 66
rect 461 38 463 66
rect 471 38 473 66
rect 481 38 483 66
rect 499 38 501 63
rect 506 38 508 63
rect 516 41 518 54
rect 529 41 531 66
rect 550 45 552 66
rect 557 45 559 66
rect 570 38 572 56
rect 598 46 600 59
rect 608 46 610 59
rect 618 39 620 57
rect 647 41 649 66
rect 660 41 662 54
rect 670 38 672 63
rect 677 38 679 63
rect 695 38 697 66
rect 705 38 707 66
rect 715 38 717 66
rect 737 38 739 66
rect 747 38 749 66
rect 757 38 759 66
rect 775 38 777 63
rect 782 38 784 63
rect 792 41 794 54
rect 805 41 807 66
rect 826 45 828 66
rect 833 45 835 66
rect 846 38 848 56
rect 874 46 876 59
rect 884 46 886 59
rect 894 39 896 57
rect 924 41 926 66
rect 937 41 939 54
rect 947 38 949 63
rect 954 38 956 63
rect 972 38 974 66
rect 982 38 984 66
rect 992 38 994 66
rect 1014 38 1016 66
rect 1024 38 1026 66
rect 1034 38 1036 66
rect 1052 38 1054 63
rect 1059 38 1061 63
rect 1069 41 1071 54
rect 1082 41 1084 66
rect 1103 45 1105 66
rect 1110 45 1112 66
rect 1123 38 1125 56
rect -149 -57 -147 -45
rect -139 -56 -137 -45
rect -129 -56 -127 -45
rect -117 -57 -115 -46
rect -97 -57 -95 -45
rect -87 -56 -85 -45
rect -77 -56 -75 -45
rect -65 -57 -63 -46
rect -45 -57 -43 -45
rect -35 -56 -33 -45
rect -25 -56 -23 -45
rect -13 -57 -11 -46
rect 7 -57 9 -45
rect 17 -56 19 -45
rect 27 -56 29 -45
rect 39 -57 41 -46
rect 59 -57 61 -45
rect 69 -56 71 -45
rect 79 -56 81 -45
rect 91 -57 93 -46
rect 112 -57 114 -45
rect 122 -56 124 -45
rect 132 -56 134 -45
rect 144 -57 146 -46
rect 169 -49 171 -37
rect 189 -49 191 -37
rect 209 -49 211 -37
rect 231 -49 233 -37
rect 253 -49 255 -37
rect 275 -49 277 -37
rect 300 -57 302 -45
rect 310 -56 312 -45
rect 320 -56 322 -45
rect 332 -57 334 -46
rect 353 -57 355 -45
rect 363 -56 365 -45
rect 373 -56 375 -45
rect 385 -57 387 -46
rect 405 -57 407 -45
rect 415 -56 417 -45
rect 425 -56 427 -45
rect 437 -57 439 -46
rect 457 -57 459 -45
rect 467 -56 469 -45
rect 477 -56 479 -45
rect 489 -57 491 -46
rect 509 -57 511 -45
rect 519 -56 521 -45
rect 529 -56 531 -45
rect 541 -57 543 -46
rect 564 -49 566 -37
rect 585 -49 587 -37
rect 608 -57 610 -45
rect 618 -56 620 -45
rect 628 -56 630 -45
rect 640 -57 642 -46
rect 661 -57 663 -45
rect 671 -56 673 -45
rect 681 -56 683 -45
rect 693 -57 695 -46
rect 713 -57 715 -45
rect 723 -56 725 -45
rect 733 -56 735 -45
rect 745 -57 747 -46
rect 765 -57 767 -45
rect 775 -56 777 -45
rect 785 -56 787 -45
rect 797 -57 799 -46
rect 817 -57 819 -45
rect 827 -56 829 -45
rect 837 -56 839 -45
rect 849 -57 851 -46
rect 869 -57 871 -45
rect 879 -56 881 -45
rect 889 -56 891 -45
rect 901 -57 903 -46
rect 922 -57 924 -45
rect 932 -56 934 -45
rect 942 -56 944 -45
rect 954 -57 956 -46
rect 976 -57 978 -45
rect 986 -56 988 -45
rect 996 -56 998 -45
rect 1008 -57 1010 -46
rect 1031 -57 1033 -45
rect 1041 -56 1043 -45
rect 1051 -56 1053 -45
rect 1063 -57 1065 -46
rect 1084 -57 1086 -45
rect 1094 -56 1096 -45
rect 1104 -56 1106 -45
rect 1116 -57 1118 -46
<< polyct0 >>
rect -244 319 -242 321
rect -234 320 -232 322
rect -200 322 -198 324
rect -206 312 -204 314
rect -150 319 -148 321
rect -140 319 -138 321
rect -118 319 -116 321
rect -108 319 -106 321
rect -58 322 -56 324
rect -11 319 -9 321
rect -52 312 -50 314
rect 32 319 34 321
rect 72 319 74 321
rect 102 322 104 324
rect 96 312 98 314
rect 152 319 154 321
rect 162 319 164 321
rect 184 319 186 321
rect 194 319 196 321
rect 244 322 246 324
rect 291 319 293 321
rect 250 312 252 314
rect 339 319 341 321
rect 379 322 381 324
rect 373 312 375 314
rect 429 319 431 321
rect 439 319 441 321
rect 461 319 463 321
rect 471 319 473 321
rect 521 322 523 324
rect 568 319 570 321
rect 527 312 529 314
rect 616 319 618 321
rect 655 322 657 324
rect 649 312 651 314
rect 705 319 707 321
rect 715 319 717 321
rect 737 319 739 321
rect 747 319 749 321
rect 797 322 799 324
rect 844 319 846 321
rect 803 312 805 314
rect 892 319 894 321
rect 932 322 934 324
rect 926 312 928 314
rect 982 319 984 321
rect 992 319 994 321
rect 1014 319 1016 321
rect 1024 319 1026 321
rect 1074 322 1076 324
rect 1121 319 1123 321
rect 1080 312 1082 314
rect -206 262 -204 264
rect -244 255 -242 257
rect -234 254 -232 256
rect -200 252 -198 254
rect -150 255 -148 257
rect -140 255 -138 257
rect -118 255 -116 257
rect -108 255 -106 257
rect -52 262 -50 264
rect -58 252 -56 254
rect -11 255 -9 257
rect 32 255 34 257
rect 72 255 74 257
rect 96 262 98 264
rect 102 252 104 254
rect 152 255 154 257
rect 162 255 164 257
rect 184 255 186 257
rect 194 255 196 257
rect 250 262 252 264
rect 244 252 246 254
rect 291 255 293 257
rect 339 255 341 257
rect 373 262 375 264
rect 379 252 381 254
rect 429 255 431 257
rect 439 255 441 257
rect 461 255 463 257
rect 471 255 473 257
rect 527 262 529 264
rect 521 252 523 254
rect 568 255 570 257
rect 616 255 618 257
rect 649 262 651 264
rect 655 252 657 254
rect 705 255 707 257
rect 715 255 717 257
rect 737 255 739 257
rect 747 255 749 257
rect 803 262 805 264
rect 797 252 799 254
rect 844 255 846 257
rect 892 255 894 257
rect 926 262 928 264
rect 932 252 934 254
rect 982 255 984 257
rect 992 255 994 257
rect 1014 255 1016 257
rect 1024 255 1026 257
rect 1080 262 1082 264
rect 1074 252 1076 254
rect 1121 255 1123 257
rect -244 175 -242 177
rect -234 176 -232 178
rect -200 178 -198 180
rect -206 168 -204 170
rect -150 175 -148 177
rect -140 175 -138 177
rect -118 175 -116 177
rect -108 175 -106 177
rect -58 178 -56 180
rect -11 175 -9 177
rect -52 168 -50 170
rect 32 175 34 177
rect 72 175 74 177
rect 102 178 104 180
rect 96 168 98 170
rect 152 175 154 177
rect 162 175 164 177
rect 184 175 186 177
rect 194 175 196 177
rect 244 178 246 180
rect 291 175 293 177
rect 250 168 252 170
rect 339 175 341 177
rect 379 178 381 180
rect 373 168 375 170
rect 429 175 431 177
rect 439 175 441 177
rect 461 175 463 177
rect 471 175 473 177
rect 521 178 523 180
rect 568 175 570 177
rect 527 168 529 170
rect 616 175 618 177
rect 655 178 657 180
rect 649 168 651 170
rect 705 175 707 177
rect 715 175 717 177
rect 737 175 739 177
rect 747 175 749 177
rect 797 178 799 180
rect 844 175 846 177
rect 803 168 805 170
rect 892 175 894 177
rect 932 178 934 180
rect 926 168 928 170
rect 982 175 984 177
rect 992 175 994 177
rect 1014 175 1016 177
rect 1024 175 1026 177
rect 1074 178 1076 180
rect 1121 175 1123 177
rect 1080 168 1082 170
rect -206 118 -204 120
rect -244 111 -242 113
rect -234 110 -232 112
rect -200 108 -198 110
rect -150 111 -148 113
rect -140 111 -138 113
rect -118 111 -116 113
rect -108 111 -106 113
rect -52 118 -50 120
rect -58 108 -56 110
rect -11 111 -9 113
rect 32 111 34 113
rect 72 111 74 113
rect 96 118 98 120
rect 102 108 104 110
rect 152 111 154 113
rect 162 111 164 113
rect 184 111 186 113
rect 194 111 196 113
rect 250 118 252 120
rect 244 108 246 110
rect 291 111 293 113
rect 339 111 341 113
rect 373 118 375 120
rect 379 108 381 110
rect 429 111 431 113
rect 439 111 441 113
rect 461 111 463 113
rect 471 111 473 113
rect 527 118 529 120
rect 521 108 523 110
rect 568 111 570 113
rect 616 111 618 113
rect 649 118 651 120
rect 655 108 657 110
rect 705 111 707 113
rect 715 111 717 113
rect 737 111 739 113
rect 747 111 749 113
rect 803 118 805 120
rect 797 108 799 110
rect 844 111 846 113
rect 892 111 894 113
rect 926 118 928 120
rect 932 108 934 110
rect 982 111 984 113
rect 992 111 994 113
rect 1014 111 1016 113
rect 1024 111 1026 113
rect 1080 118 1082 120
rect 1074 108 1076 110
rect 1121 111 1123 113
rect -244 31 -242 33
rect -234 32 -232 34
rect -200 34 -198 36
rect -206 24 -204 26
rect -150 31 -148 33
rect -140 31 -138 33
rect -118 31 -116 33
rect -108 31 -106 33
rect -58 34 -56 36
rect -11 31 -9 33
rect -52 24 -50 26
rect 32 31 34 33
rect 72 31 74 33
rect 102 34 104 36
rect 96 24 98 26
rect 152 31 154 33
rect 162 31 164 33
rect 184 31 186 33
rect 194 31 196 33
rect 244 34 246 36
rect 291 31 293 33
rect 250 24 252 26
rect 339 31 341 33
rect 379 34 381 36
rect 373 24 375 26
rect 429 31 431 33
rect 439 31 441 33
rect 461 31 463 33
rect 471 31 473 33
rect 521 34 523 36
rect 568 31 570 33
rect 527 24 529 26
rect 616 31 618 33
rect 655 34 657 36
rect 649 24 651 26
rect 705 31 707 33
rect 715 31 717 33
rect 737 31 739 33
rect 747 31 749 33
rect 797 34 799 36
rect 844 31 846 33
rect 803 24 805 26
rect 892 31 894 33
rect 932 34 934 36
rect 926 24 928 26
rect 982 31 984 33
rect 992 31 994 33
rect 1014 31 1016 33
rect 1024 31 1026 33
rect 1074 34 1076 36
rect 1121 31 1123 33
rect 1080 24 1082 26
rect -147 -33 -145 -31
rect -95 -33 -93 -31
rect -43 -33 -41 -31
rect 9 -33 11 -31
rect 61 -33 63 -31
rect 114 -33 116 -31
rect 302 -33 304 -31
rect 355 -33 357 -31
rect 407 -33 409 -31
rect 459 -33 461 -31
rect 511 -33 513 -31
rect 610 -33 612 -31
rect 663 -33 665 -31
rect 715 -33 717 -31
rect 767 -33 769 -31
rect 819 -33 821 -31
rect 871 -33 873 -31
rect 924 -33 926 -31
rect 978 -33 980 -31
rect 1033 -33 1035 -31
rect 1086 -33 1088 -31
<< polyct1 >>
rect -281 327 -279 329
rect -265 314 -263 316
rect -186 319 -184 321
rect -167 319 -165 321
rect -160 319 -158 321
rect -98 319 -96 321
rect -91 319 -89 321
rect -72 319 -70 321
rect -31 326 -29 328
rect 12 327 14 329
rect -21 319 -19 321
rect 52 327 54 329
rect 22 319 24 321
rect 62 319 64 321
rect 116 319 118 321
rect 135 319 137 321
rect 142 319 144 321
rect 204 319 206 321
rect 211 319 213 321
rect 230 319 232 321
rect 271 326 273 328
rect 319 327 321 329
rect 281 319 283 321
rect 329 319 331 321
rect 393 319 395 321
rect 412 319 414 321
rect 419 319 421 321
rect 481 319 483 321
rect 488 319 490 321
rect 507 319 509 321
rect 548 326 550 328
rect 596 327 598 329
rect 558 319 560 321
rect 606 319 608 321
rect 669 319 671 321
rect 688 319 690 321
rect 695 319 697 321
rect 757 319 759 321
rect 764 319 766 321
rect 783 319 785 321
rect 824 326 826 328
rect 872 327 874 329
rect 834 319 836 321
rect 882 319 884 321
rect 946 319 948 321
rect 965 319 967 321
rect 972 319 974 321
rect 1034 319 1036 321
rect 1041 319 1043 321
rect 1060 319 1062 321
rect 1101 326 1103 328
rect 1111 319 1113 321
rect -265 260 -263 262
rect -281 247 -279 249
rect -186 255 -184 257
rect -167 255 -165 257
rect -160 255 -158 257
rect -98 255 -96 257
rect -91 255 -89 257
rect -72 255 -70 257
rect -21 255 -19 257
rect -31 248 -29 250
rect 22 255 24 257
rect 12 247 14 249
rect 62 255 64 257
rect 52 247 54 249
rect 116 255 118 257
rect 135 255 137 257
rect 142 255 144 257
rect 204 255 206 257
rect 211 255 213 257
rect 230 255 232 257
rect 281 255 283 257
rect 271 248 273 250
rect 329 255 331 257
rect 319 247 321 249
rect 393 255 395 257
rect 412 255 414 257
rect 419 255 421 257
rect 481 255 483 257
rect 488 255 490 257
rect 507 255 509 257
rect 558 255 560 257
rect 548 248 550 250
rect 606 255 608 257
rect 596 247 598 249
rect 669 255 671 257
rect 688 255 690 257
rect 695 255 697 257
rect 757 255 759 257
rect 764 255 766 257
rect 783 255 785 257
rect 834 255 836 257
rect 824 248 826 250
rect 882 255 884 257
rect 872 247 874 249
rect 946 255 948 257
rect 965 255 967 257
rect 972 255 974 257
rect 1034 255 1036 257
rect 1041 255 1043 257
rect 1060 255 1062 257
rect 1111 255 1113 257
rect 1101 248 1103 250
rect -281 183 -279 185
rect -265 170 -263 172
rect -186 175 -184 177
rect -167 175 -165 177
rect -160 175 -158 177
rect -98 175 -96 177
rect -91 175 -89 177
rect -72 175 -70 177
rect -31 182 -29 184
rect 12 183 14 185
rect -21 175 -19 177
rect 52 183 54 185
rect 22 175 24 177
rect 62 175 64 177
rect 116 175 118 177
rect 135 175 137 177
rect 142 175 144 177
rect 204 175 206 177
rect 211 175 213 177
rect 230 175 232 177
rect 271 182 273 184
rect 319 183 321 185
rect 281 175 283 177
rect 329 175 331 177
rect 393 175 395 177
rect 412 175 414 177
rect 419 175 421 177
rect 481 175 483 177
rect 488 175 490 177
rect 507 175 509 177
rect 548 182 550 184
rect 596 183 598 185
rect 558 175 560 177
rect 606 175 608 177
rect 669 175 671 177
rect 688 175 690 177
rect 695 175 697 177
rect 757 175 759 177
rect 764 175 766 177
rect 783 175 785 177
rect 824 182 826 184
rect 872 183 874 185
rect 834 175 836 177
rect 882 175 884 177
rect 946 175 948 177
rect 965 175 967 177
rect 972 175 974 177
rect 1034 175 1036 177
rect 1041 175 1043 177
rect 1060 175 1062 177
rect 1101 182 1103 184
rect 1111 175 1113 177
rect -265 116 -263 118
rect -281 103 -279 105
rect -186 111 -184 113
rect -167 111 -165 113
rect -160 111 -158 113
rect -98 111 -96 113
rect -91 111 -89 113
rect -72 111 -70 113
rect -21 111 -19 113
rect -31 104 -29 106
rect 22 111 24 113
rect 12 103 14 105
rect 62 111 64 113
rect 52 103 54 105
rect 116 111 118 113
rect 135 111 137 113
rect 142 111 144 113
rect 204 111 206 113
rect 211 111 213 113
rect 230 111 232 113
rect 281 111 283 113
rect 271 104 273 106
rect 329 111 331 113
rect 319 103 321 105
rect 393 111 395 113
rect 412 111 414 113
rect 419 111 421 113
rect 481 111 483 113
rect 488 111 490 113
rect 507 111 509 113
rect 558 111 560 113
rect 548 104 550 106
rect 606 111 608 113
rect 596 103 598 105
rect 669 111 671 113
rect 688 111 690 113
rect 695 111 697 113
rect 757 111 759 113
rect 764 111 766 113
rect 783 111 785 113
rect 834 111 836 113
rect 824 104 826 106
rect 882 111 884 113
rect 872 103 874 105
rect 946 111 948 113
rect 965 111 967 113
rect 972 111 974 113
rect 1034 111 1036 113
rect 1041 111 1043 113
rect 1060 111 1062 113
rect 1111 111 1113 113
rect 1101 104 1103 106
rect -281 39 -279 41
rect -265 26 -263 28
rect -186 31 -184 33
rect -167 31 -165 33
rect -160 31 -158 33
rect -98 31 -96 33
rect -91 31 -89 33
rect -72 31 -70 33
rect -31 38 -29 40
rect 12 39 14 41
rect -21 31 -19 33
rect 52 39 54 41
rect 22 31 24 33
rect 62 31 64 33
rect 116 31 118 33
rect 135 31 137 33
rect 142 31 144 33
rect 204 31 206 33
rect 211 31 213 33
rect 230 31 232 33
rect 271 38 273 40
rect 319 39 321 41
rect 281 31 283 33
rect 329 31 331 33
rect 393 31 395 33
rect 412 31 414 33
rect 419 31 421 33
rect 481 31 483 33
rect 488 31 490 33
rect 507 31 509 33
rect 548 38 550 40
rect 596 39 598 41
rect 558 31 560 33
rect 606 31 608 33
rect 669 31 671 33
rect 688 31 690 33
rect 695 31 697 33
rect 757 31 759 33
rect 764 31 766 33
rect 783 31 785 33
rect 824 38 826 40
rect 872 39 874 41
rect 834 31 836 33
rect 882 31 884 33
rect 946 31 948 33
rect 965 31 967 33
rect 972 31 974 33
rect 1034 31 1036 33
rect 1041 31 1043 33
rect 1060 31 1062 33
rect 1101 38 1103 40
rect 1111 31 1113 33
rect -137 -32 -135 -30
rect -115 -32 -113 -30
rect -125 -40 -123 -38
rect -85 -32 -83 -30
rect -63 -32 -61 -30
rect -73 -40 -71 -38
rect -33 -32 -31 -30
rect -11 -32 -9 -30
rect -21 -40 -19 -38
rect 19 -32 21 -30
rect 41 -32 43 -30
rect 31 -40 33 -38
rect 71 -32 73 -30
rect 93 -32 95 -30
rect 83 -40 85 -38
rect 124 -32 126 -30
rect 146 -32 148 -30
rect 136 -40 138 -38
rect 312 -32 314 -30
rect 334 -32 336 -30
rect 324 -40 326 -38
rect 171 -56 173 -54
rect 191 -56 193 -54
rect 211 -56 213 -54
rect 233 -56 235 -54
rect 255 -56 257 -54
rect 277 -56 279 -54
rect 365 -32 367 -30
rect 387 -32 389 -30
rect 377 -40 379 -38
rect 417 -32 419 -30
rect 439 -32 441 -30
rect 429 -40 431 -38
rect 469 -32 471 -30
rect 491 -32 493 -30
rect 481 -40 483 -38
rect 521 -32 523 -30
rect 543 -32 545 -30
rect 533 -40 535 -38
rect 620 -32 622 -30
rect 642 -32 644 -30
rect 632 -40 634 -38
rect 566 -56 568 -54
rect 587 -56 589 -54
rect 673 -32 675 -30
rect 695 -32 697 -30
rect 685 -40 687 -38
rect 725 -32 727 -30
rect 747 -32 749 -30
rect 737 -40 739 -38
rect 777 -32 779 -30
rect 799 -32 801 -30
rect 789 -40 791 -38
rect 829 -32 831 -30
rect 851 -32 853 -30
rect 841 -40 843 -38
rect 881 -32 883 -30
rect 903 -32 905 -30
rect 893 -40 895 -38
rect 934 -32 936 -30
rect 956 -32 958 -30
rect 946 -40 948 -38
rect 988 -32 990 -30
rect 1010 -32 1012 -30
rect 1000 -40 1002 -38
rect 1043 -32 1045 -30
rect 1065 -32 1067 -30
rect 1055 -40 1057 -38
rect 1096 -32 1098 -30
rect 1118 -32 1120 -30
rect 1108 -40 1110 -38
<< ndifct0 >>
rect -281 310 -279 312
rect -267 302 -265 304
rect -255 305 -253 307
rect -203 299 -201 301
rect -193 302 -191 304
rect -183 310 -181 312
rect -173 310 -171 312
rect -173 303 -171 305
rect -163 303 -161 305
rect -146 296 -144 298
rect -112 296 -110 298
rect -85 310 -83 312
rect -95 303 -93 305
rect -85 303 -83 305
rect -75 310 -73 312
rect -24 310 -22 312
rect -65 302 -63 304
rect -55 299 -53 301
rect -34 297 -32 299
rect 9 303 11 305
rect 49 303 51 305
rect -15 297 -13 299
rect 99 299 101 301
rect 109 302 111 304
rect 119 310 121 312
rect 129 310 131 312
rect 129 303 131 305
rect 139 303 141 305
rect 156 296 158 298
rect 190 296 192 298
rect 217 310 219 312
rect 207 303 209 305
rect 217 303 219 305
rect 227 310 229 312
rect 278 310 280 312
rect 237 302 239 304
rect 247 299 249 301
rect 268 297 270 299
rect 316 303 318 305
rect 287 297 289 299
rect 376 299 378 301
rect 386 302 388 304
rect 396 310 398 312
rect 406 310 408 312
rect 406 303 408 305
rect 416 303 418 305
rect 433 296 435 298
rect 467 296 469 298
rect 494 310 496 312
rect 484 303 486 305
rect 494 303 496 305
rect 504 310 506 312
rect 555 310 557 312
rect 514 302 516 304
rect 524 299 526 301
rect 545 297 547 299
rect 593 303 595 305
rect 564 297 566 299
rect 652 299 654 301
rect 662 302 664 304
rect 672 310 674 312
rect 682 310 684 312
rect 682 303 684 305
rect 692 303 694 305
rect 709 296 711 298
rect 743 296 745 298
rect 770 310 772 312
rect 760 303 762 305
rect 770 303 772 305
rect 780 310 782 312
rect 831 310 833 312
rect 790 302 792 304
rect 800 299 802 301
rect 821 297 823 299
rect 869 303 871 305
rect 840 297 842 299
rect 929 299 931 301
rect 939 302 941 304
rect 949 310 951 312
rect 959 310 961 312
rect 959 303 961 305
rect 969 303 971 305
rect 986 296 988 298
rect 1020 296 1022 298
rect 1047 310 1049 312
rect 1037 303 1039 305
rect 1047 303 1049 305
rect 1057 310 1059 312
rect 1108 310 1110 312
rect 1067 302 1069 304
rect 1077 299 1079 301
rect 1098 297 1100 299
rect 1117 297 1119 299
rect -267 272 -265 274
rect -281 264 -279 266
rect -255 269 -253 271
rect -203 275 -201 277
rect -193 272 -191 274
rect -183 264 -181 266
rect -173 271 -171 273
rect -163 271 -161 273
rect -173 264 -171 266
rect -146 278 -144 280
rect -112 278 -110 280
rect -95 271 -93 273
rect -85 271 -83 273
rect -85 264 -83 266
rect -75 264 -73 266
rect -65 272 -63 274
rect -55 275 -53 277
rect -34 277 -32 279
rect -15 277 -13 279
rect 9 271 11 273
rect -24 264 -22 266
rect 49 271 51 273
rect 99 275 101 277
rect 109 272 111 274
rect 119 264 121 266
rect 129 271 131 273
rect 139 271 141 273
rect 129 264 131 266
rect 156 278 158 280
rect 190 278 192 280
rect 207 271 209 273
rect 217 271 219 273
rect 217 264 219 266
rect 227 264 229 266
rect 237 272 239 274
rect 247 275 249 277
rect 268 277 270 279
rect 287 277 289 279
rect 316 271 318 273
rect 278 264 280 266
rect 376 275 378 277
rect 386 272 388 274
rect 396 264 398 266
rect 406 271 408 273
rect 416 271 418 273
rect 406 264 408 266
rect 433 278 435 280
rect 467 278 469 280
rect 484 271 486 273
rect 494 271 496 273
rect 494 264 496 266
rect 504 264 506 266
rect 514 272 516 274
rect 524 275 526 277
rect 545 277 547 279
rect 564 277 566 279
rect 593 271 595 273
rect 555 264 557 266
rect 652 275 654 277
rect 662 272 664 274
rect 672 264 674 266
rect 682 271 684 273
rect 692 271 694 273
rect 682 264 684 266
rect 709 278 711 280
rect 743 278 745 280
rect 760 271 762 273
rect 770 271 772 273
rect 770 264 772 266
rect 780 264 782 266
rect 790 272 792 274
rect 800 275 802 277
rect 821 277 823 279
rect 840 277 842 279
rect 869 271 871 273
rect 831 264 833 266
rect 929 275 931 277
rect 939 272 941 274
rect 949 264 951 266
rect 959 271 961 273
rect 969 271 971 273
rect 959 264 961 266
rect 986 278 988 280
rect 1020 278 1022 280
rect 1037 271 1039 273
rect 1047 271 1049 273
rect 1047 264 1049 266
rect 1057 264 1059 266
rect 1067 272 1069 274
rect 1077 275 1079 277
rect 1098 277 1100 279
rect 1117 277 1119 279
rect 1108 264 1110 266
rect -281 166 -279 168
rect -267 158 -265 160
rect -255 161 -253 163
rect -203 155 -201 157
rect -193 158 -191 160
rect -183 166 -181 168
rect -173 166 -171 168
rect -173 159 -171 161
rect -163 159 -161 161
rect -146 152 -144 154
rect -112 152 -110 154
rect -85 166 -83 168
rect -95 159 -93 161
rect -85 159 -83 161
rect -75 166 -73 168
rect -24 166 -22 168
rect -65 158 -63 160
rect -55 155 -53 157
rect -34 153 -32 155
rect 9 159 11 161
rect 49 159 51 161
rect -15 153 -13 155
rect 99 155 101 157
rect 109 158 111 160
rect 119 166 121 168
rect 129 166 131 168
rect 129 159 131 161
rect 139 159 141 161
rect 156 152 158 154
rect 190 152 192 154
rect 217 166 219 168
rect 207 159 209 161
rect 217 159 219 161
rect 227 166 229 168
rect 278 166 280 168
rect 237 158 239 160
rect 247 155 249 157
rect 268 153 270 155
rect 316 159 318 161
rect 287 153 289 155
rect 376 155 378 157
rect 386 158 388 160
rect 396 166 398 168
rect 406 166 408 168
rect 406 159 408 161
rect 416 159 418 161
rect 433 152 435 154
rect 467 152 469 154
rect 494 166 496 168
rect 484 159 486 161
rect 494 159 496 161
rect 504 166 506 168
rect 555 166 557 168
rect 514 158 516 160
rect 524 155 526 157
rect 545 153 547 155
rect 593 159 595 161
rect 564 153 566 155
rect 652 155 654 157
rect 662 158 664 160
rect 672 166 674 168
rect 682 166 684 168
rect 682 159 684 161
rect 692 159 694 161
rect 709 152 711 154
rect 743 152 745 154
rect 770 166 772 168
rect 760 159 762 161
rect 770 159 772 161
rect 780 166 782 168
rect 831 166 833 168
rect 790 158 792 160
rect 800 155 802 157
rect 821 153 823 155
rect 869 159 871 161
rect 840 153 842 155
rect 929 155 931 157
rect 939 158 941 160
rect 949 166 951 168
rect 959 166 961 168
rect 959 159 961 161
rect 969 159 971 161
rect 986 152 988 154
rect 1020 152 1022 154
rect 1047 166 1049 168
rect 1037 159 1039 161
rect 1047 159 1049 161
rect 1057 166 1059 168
rect 1108 166 1110 168
rect 1067 158 1069 160
rect 1077 155 1079 157
rect 1098 153 1100 155
rect 1117 153 1119 155
rect -267 128 -265 130
rect -281 120 -279 122
rect -255 125 -253 127
rect -203 131 -201 133
rect -193 128 -191 130
rect -183 120 -181 122
rect -173 127 -171 129
rect -163 127 -161 129
rect -173 120 -171 122
rect -146 134 -144 136
rect -112 134 -110 136
rect -95 127 -93 129
rect -85 127 -83 129
rect -85 120 -83 122
rect -75 120 -73 122
rect -65 128 -63 130
rect -55 131 -53 133
rect -34 133 -32 135
rect -15 133 -13 135
rect 9 127 11 129
rect -24 120 -22 122
rect 49 127 51 129
rect 99 131 101 133
rect 109 128 111 130
rect 119 120 121 122
rect 129 127 131 129
rect 139 127 141 129
rect 129 120 131 122
rect 156 134 158 136
rect 190 134 192 136
rect 207 127 209 129
rect 217 127 219 129
rect 217 120 219 122
rect 227 120 229 122
rect 237 128 239 130
rect 247 131 249 133
rect 268 133 270 135
rect 287 133 289 135
rect 316 127 318 129
rect 278 120 280 122
rect 376 131 378 133
rect 386 128 388 130
rect 396 120 398 122
rect 406 127 408 129
rect 416 127 418 129
rect 406 120 408 122
rect 433 134 435 136
rect 467 134 469 136
rect 484 127 486 129
rect 494 127 496 129
rect 494 120 496 122
rect 504 120 506 122
rect 514 128 516 130
rect 524 131 526 133
rect 545 133 547 135
rect 564 133 566 135
rect 593 127 595 129
rect 555 120 557 122
rect 652 131 654 133
rect 662 128 664 130
rect 672 120 674 122
rect 682 127 684 129
rect 692 127 694 129
rect 682 120 684 122
rect 709 134 711 136
rect 743 134 745 136
rect 760 127 762 129
rect 770 127 772 129
rect 770 120 772 122
rect 780 120 782 122
rect 790 128 792 130
rect 800 131 802 133
rect 821 133 823 135
rect 840 133 842 135
rect 869 127 871 129
rect 831 120 833 122
rect 929 131 931 133
rect 939 128 941 130
rect 949 120 951 122
rect 959 127 961 129
rect 969 127 971 129
rect 959 120 961 122
rect 986 134 988 136
rect 1020 134 1022 136
rect 1037 127 1039 129
rect 1047 127 1049 129
rect 1047 120 1049 122
rect 1057 120 1059 122
rect 1067 128 1069 130
rect 1077 131 1079 133
rect 1098 133 1100 135
rect 1117 133 1119 135
rect 1108 120 1110 122
rect -281 22 -279 24
rect -267 14 -265 16
rect -255 17 -253 19
rect -203 11 -201 13
rect -193 14 -191 16
rect -183 22 -181 24
rect -173 22 -171 24
rect -173 15 -171 17
rect -163 15 -161 17
rect -146 8 -144 10
rect -112 8 -110 10
rect -85 22 -83 24
rect -95 15 -93 17
rect -85 15 -83 17
rect -75 22 -73 24
rect -24 22 -22 24
rect -65 14 -63 16
rect -55 11 -53 13
rect -34 9 -32 11
rect 9 15 11 17
rect 49 15 51 17
rect -15 9 -13 11
rect 99 11 101 13
rect 109 14 111 16
rect 119 22 121 24
rect 129 22 131 24
rect 129 15 131 17
rect 139 15 141 17
rect 156 8 158 10
rect 190 8 192 10
rect 217 22 219 24
rect 207 15 209 17
rect 217 15 219 17
rect 227 22 229 24
rect 278 22 280 24
rect 237 14 239 16
rect 247 11 249 13
rect 268 9 270 11
rect 316 15 318 17
rect 287 9 289 11
rect 376 11 378 13
rect 386 14 388 16
rect 396 22 398 24
rect 406 22 408 24
rect 406 15 408 17
rect 416 15 418 17
rect 433 8 435 10
rect 467 8 469 10
rect 494 22 496 24
rect 484 15 486 17
rect 494 15 496 17
rect 504 22 506 24
rect 555 22 557 24
rect 514 14 516 16
rect 524 11 526 13
rect 545 9 547 11
rect 593 15 595 17
rect 564 9 566 11
rect 652 11 654 13
rect 662 14 664 16
rect 672 22 674 24
rect 682 22 684 24
rect 682 15 684 17
rect 692 15 694 17
rect 709 8 711 10
rect 743 8 745 10
rect 770 22 772 24
rect 760 15 762 17
rect 770 15 772 17
rect 780 22 782 24
rect 831 22 833 24
rect 790 14 792 16
rect 800 11 802 13
rect 821 9 823 11
rect 869 15 871 17
rect 840 9 842 11
rect 929 11 931 13
rect 939 14 941 16
rect 949 22 951 24
rect 959 22 961 24
rect 959 15 961 17
rect 969 15 971 17
rect 986 8 988 10
rect 1020 8 1022 10
rect 1047 22 1049 24
rect 1037 15 1039 17
rect 1047 15 1049 17
rect 1057 22 1059 24
rect 1108 22 1110 24
rect 1067 14 1069 16
rect 1077 11 1079 13
rect 1098 9 1100 11
rect 1117 9 1119 11
rect -115 -18 -113 -16
rect -63 -18 -61 -16
rect -11 -18 -9 -16
rect 41 -18 43 -16
rect 93 -18 95 -16
rect 146 -18 148 -16
rect 174 -23 176 -21
rect 194 -23 196 -21
rect 214 -23 216 -21
rect 236 -23 238 -21
rect 258 -23 260 -21
rect 280 -23 282 -21
rect 334 -18 336 -16
rect 387 -18 389 -16
rect 439 -18 441 -16
rect 491 -18 493 -16
rect 543 -18 545 -16
rect 569 -23 571 -21
rect 590 -23 592 -21
rect 642 -18 644 -16
rect 695 -18 697 -16
rect 747 -18 749 -16
rect 799 -18 801 -16
rect 851 -18 853 -16
rect 903 -18 905 -16
rect 956 -18 958 -16
rect 1010 -18 1012 -16
rect 1065 -18 1067 -16
rect 1118 -18 1120 -16
<< ndifct1 >>
rect -245 303 -243 305
rect -213 303 -211 305
rect -227 293 -225 295
rect -135 303 -133 305
rect -123 303 -121 305
rect -45 303 -43 305
rect -4 310 -2 312
rect 39 305 41 307
rect 79 305 81 307
rect 89 303 91 305
rect 28 293 30 295
rect 68 293 70 295
rect 167 303 169 305
rect 179 303 181 305
rect 257 303 259 305
rect 298 310 300 312
rect 346 305 348 307
rect 366 303 368 305
rect 335 293 337 295
rect 444 303 446 305
rect 456 303 458 305
rect 534 303 536 305
rect 575 310 577 312
rect 623 305 625 307
rect 642 303 644 305
rect 612 293 614 295
rect 720 303 722 305
rect 732 303 734 305
rect 810 303 812 305
rect 851 310 853 312
rect 899 305 901 307
rect 919 303 921 305
rect 888 293 890 295
rect 997 303 999 305
rect 1009 303 1011 305
rect 1087 303 1089 305
rect 1128 310 1130 312
rect -227 281 -225 283
rect -245 271 -243 273
rect -213 271 -211 273
rect -135 271 -133 273
rect -123 271 -121 273
rect 28 281 30 283
rect -45 271 -43 273
rect 68 281 70 283
rect -4 264 -2 266
rect 39 269 41 271
rect 79 269 81 271
rect 89 271 91 273
rect 167 271 169 273
rect 179 271 181 273
rect 335 281 337 283
rect 257 271 259 273
rect 298 264 300 266
rect 346 269 348 271
rect 366 271 368 273
rect 444 271 446 273
rect 456 271 458 273
rect 612 281 614 283
rect 534 271 536 273
rect 575 264 577 266
rect 623 269 625 271
rect 642 271 644 273
rect 720 271 722 273
rect 732 271 734 273
rect 888 281 890 283
rect 810 271 812 273
rect 851 264 853 266
rect 899 269 901 271
rect 919 271 921 273
rect 997 271 999 273
rect 1009 271 1011 273
rect 1087 271 1089 273
rect 1128 264 1130 266
rect -245 159 -243 161
rect -213 159 -211 161
rect -227 149 -225 151
rect -135 159 -133 161
rect -123 159 -121 161
rect -45 159 -43 161
rect -4 166 -2 168
rect 39 161 41 163
rect 79 161 81 163
rect 89 159 91 161
rect 28 149 30 151
rect 68 149 70 151
rect 167 159 169 161
rect 179 159 181 161
rect 257 159 259 161
rect 298 166 300 168
rect 346 161 348 163
rect 366 159 368 161
rect 335 149 337 151
rect 444 159 446 161
rect 456 159 458 161
rect 534 159 536 161
rect 575 166 577 168
rect 623 161 625 163
rect 642 159 644 161
rect 612 149 614 151
rect 720 159 722 161
rect 732 159 734 161
rect 810 159 812 161
rect 851 166 853 168
rect 899 161 901 163
rect 919 159 921 161
rect 888 149 890 151
rect 997 159 999 161
rect 1009 159 1011 161
rect 1087 159 1089 161
rect 1128 166 1130 168
rect -227 137 -225 139
rect -245 127 -243 129
rect -213 127 -211 129
rect -135 127 -133 129
rect -123 127 -121 129
rect 28 137 30 139
rect -45 127 -43 129
rect 68 137 70 139
rect -4 120 -2 122
rect 39 125 41 127
rect 79 125 81 127
rect 89 127 91 129
rect 167 127 169 129
rect 179 127 181 129
rect 335 137 337 139
rect 257 127 259 129
rect 298 120 300 122
rect 346 125 348 127
rect 366 127 368 129
rect 444 127 446 129
rect 456 127 458 129
rect 612 137 614 139
rect 534 127 536 129
rect 575 120 577 122
rect 623 125 625 127
rect 642 127 644 129
rect 720 127 722 129
rect 732 127 734 129
rect 888 137 890 139
rect 810 127 812 129
rect 851 120 853 122
rect 899 125 901 127
rect 919 127 921 129
rect 997 127 999 129
rect 1009 127 1011 129
rect 1087 127 1089 129
rect 1128 120 1130 122
rect -245 15 -243 17
rect -213 15 -211 17
rect -227 5 -225 7
rect -135 15 -133 17
rect -123 15 -121 17
rect -45 15 -43 17
rect -4 22 -2 24
rect 39 17 41 19
rect 79 17 81 19
rect 89 15 91 17
rect 28 5 30 7
rect 68 5 70 7
rect 167 15 169 17
rect 179 15 181 17
rect 257 15 259 17
rect 298 22 300 24
rect 346 17 348 19
rect 366 15 368 17
rect 335 5 337 7
rect 444 15 446 17
rect 456 15 458 17
rect 534 15 536 17
rect 575 22 577 24
rect 623 17 625 19
rect 642 15 644 17
rect 612 5 614 7
rect 720 15 722 17
rect 732 15 734 17
rect 810 15 812 17
rect 851 22 853 24
rect 899 17 901 19
rect 919 15 921 17
rect 888 5 890 7
rect 997 15 999 17
rect 1009 15 1011 17
rect 1087 15 1089 17
rect 1128 22 1130 24
rect -142 -6 -140 -4
rect -90 -6 -88 -4
rect -38 -6 -36 -4
rect 14 -6 16 -4
rect 66 -6 68 -4
rect 119 -6 121 -4
rect 307 -6 309 -4
rect 360 -6 362 -4
rect 412 -6 414 -4
rect 464 -6 466 -4
rect 516 -6 518 -4
rect 615 -6 617 -4
rect 668 -6 670 -4
rect 720 -6 722 -4
rect 772 -6 774 -4
rect 824 -6 826 -4
rect 876 -6 878 -4
rect 929 -6 931 -4
rect 983 -6 985 -4
rect 1038 -6 1040 -4
rect 1091 -6 1093 -4
rect -154 -23 -152 -21
rect -102 -23 -100 -21
rect -50 -23 -48 -21
rect 2 -23 4 -21
rect 54 -23 56 -21
rect 107 -23 109 -21
rect 164 -23 166 -21
rect 184 -23 186 -21
rect 204 -23 206 -21
rect 226 -23 228 -21
rect 248 -23 250 -21
rect 270 -23 272 -21
rect 295 -23 297 -21
rect 348 -23 350 -21
rect 400 -23 402 -21
rect 452 -23 454 -21
rect 504 -23 506 -21
rect 559 -23 561 -21
rect 580 -23 582 -21
rect 603 -23 605 -21
rect 656 -23 658 -21
rect 708 -23 710 -21
rect 760 -23 762 -21
rect 812 -23 814 -21
rect 864 -23 866 -21
rect 917 -23 919 -21
rect 971 -23 973 -21
rect 1026 -23 1028 -21
rect 1079 -23 1081 -21
<< ntiect1 >>
rect -247 353 -245 355
rect -5 353 -3 355
rect 38 353 40 355
rect 78 353 80 355
rect 297 353 299 355
rect 345 353 347 355
rect 574 353 576 355
rect 622 353 624 355
rect 850 353 852 355
rect 898 353 900 355
rect 1127 353 1129 355
rect -247 221 -245 223
rect -5 221 -3 223
rect 38 221 40 223
rect 78 221 80 223
rect 297 221 299 223
rect 345 221 347 223
rect 574 221 576 223
rect 622 221 624 223
rect 850 221 852 223
rect 898 221 900 223
rect 1127 221 1129 223
rect -247 209 -245 211
rect -5 209 -3 211
rect 38 209 40 211
rect 78 209 80 211
rect 297 209 299 211
rect 345 209 347 211
rect 574 209 576 211
rect 622 209 624 211
rect 850 209 852 211
rect 898 209 900 211
rect 1127 209 1129 211
rect -247 77 -245 79
rect -5 77 -3 79
rect 38 77 40 79
rect 78 77 80 79
rect 297 77 299 79
rect 345 77 347 79
rect 574 77 576 79
rect 622 77 624 79
rect 850 77 852 79
rect 898 77 900 79
rect 1127 77 1129 79
rect -247 65 -245 67
rect -5 65 -3 67
rect 38 65 40 67
rect 78 65 80 67
rect 297 65 299 67
rect 345 65 347 67
rect 574 65 576 67
rect 622 65 624 67
rect 850 65 852 67
rect 898 65 900 67
rect 1127 65 1129 67
rect -133 -66 -131 -64
rect -81 -66 -79 -64
rect -29 -66 -27 -64
rect 23 -66 25 -64
rect 75 -66 77 -64
rect 128 -66 130 -64
rect 174 -66 176 -64
rect 194 -66 196 -64
rect 214 -66 216 -64
rect 236 -66 238 -64
rect 258 -66 260 -64
rect 280 -66 282 -64
rect 316 -66 318 -64
rect 369 -66 371 -64
rect 421 -66 423 -64
rect 473 -66 475 -64
rect 525 -66 527 -64
rect 569 -66 571 -64
rect 590 -66 592 -64
rect 624 -66 626 -64
rect 677 -66 679 -64
rect 729 -66 731 -64
rect 781 -66 783 -64
rect 833 -66 835 -64
rect 885 -66 887 -64
rect 938 -66 940 -64
rect 992 -66 994 -64
rect 1047 -66 1049 -64
rect 1100 -66 1102 -64
<< ptiect1 >>
rect -280 293 -278 295
rect -5 293 -3 295
rect 38 293 40 295
rect 78 293 80 295
rect 297 293 299 295
rect 345 293 347 295
rect 574 293 576 295
rect 622 293 624 295
rect 850 293 852 295
rect 898 293 900 295
rect 1127 293 1129 295
rect -280 281 -278 283
rect -5 281 -3 283
rect 38 281 40 283
rect 78 281 80 283
rect 297 281 299 283
rect 345 281 347 283
rect 574 281 576 283
rect 622 281 624 283
rect 850 281 852 283
rect 898 281 900 283
rect 1127 281 1129 283
rect -280 149 -278 151
rect -5 149 -3 151
rect 38 149 40 151
rect 78 149 80 151
rect 297 149 299 151
rect 345 149 347 151
rect 574 149 576 151
rect 622 149 624 151
rect 850 149 852 151
rect 898 149 900 151
rect 1127 149 1129 151
rect -280 137 -278 139
rect -5 137 -3 139
rect 38 137 40 139
rect 78 137 80 139
rect 297 137 299 139
rect 345 137 347 139
rect 574 137 576 139
rect 622 137 624 139
rect 850 137 852 139
rect 898 137 900 139
rect 1127 137 1129 139
rect -280 5 -278 7
rect -5 5 -3 7
rect 38 5 40 7
rect 78 5 80 7
rect 297 5 299 7
rect 345 5 347 7
rect 574 5 576 7
rect 622 5 624 7
rect 850 5 852 7
rect 898 5 900 7
rect 1127 5 1129 7
rect -153 -6 -151 -4
rect -121 -6 -119 -4
rect -113 -6 -111 -4
rect -101 -6 -99 -4
rect -69 -6 -67 -4
rect -61 -6 -59 -4
rect -49 -6 -47 -4
rect -17 -6 -15 -4
rect -9 -6 -7 -4
rect 3 -6 5 -4
rect 35 -6 37 -4
rect 43 -6 45 -4
rect 55 -6 57 -4
rect 87 -6 89 -4
rect 95 -6 97 -4
rect 108 -6 110 -4
rect 140 -6 142 -4
rect 148 -6 150 -4
rect 165 -6 167 -4
rect 173 -6 175 -4
rect 185 -6 187 -4
rect 193 -6 195 -4
rect 205 -6 207 -4
rect 213 -6 215 -4
rect 227 -6 229 -4
rect 235 -6 237 -4
rect 249 -6 251 -4
rect 257 -6 259 -4
rect 271 -6 273 -4
rect 279 -6 281 -4
rect 296 -6 298 -4
rect 328 -6 330 -4
rect 336 -6 338 -4
rect 349 -6 351 -4
rect 381 -6 383 -4
rect 389 -6 391 -4
rect 401 -6 403 -4
rect 433 -6 435 -4
rect 441 -6 443 -4
rect 453 -6 455 -4
rect 485 -6 487 -4
rect 493 -6 495 -4
rect 505 -6 507 -4
rect 537 -6 539 -4
rect 545 -6 547 -4
rect 560 -6 562 -4
rect 568 -6 570 -4
rect 581 -6 583 -4
rect 589 -6 591 -4
rect 604 -6 606 -4
rect 636 -6 638 -4
rect 644 -6 646 -4
rect 657 -6 659 -4
rect 689 -6 691 -4
rect 697 -6 699 -4
rect 709 -6 711 -4
rect 741 -6 743 -4
rect 749 -6 751 -4
rect 761 -6 763 -4
rect 793 -6 795 -4
rect 801 -6 803 -4
rect 813 -6 815 -4
rect 845 -6 847 -4
rect 853 -6 855 -4
rect 865 -6 867 -4
rect 897 -6 899 -4
rect 905 -6 907 -4
rect 918 -6 920 -4
rect 950 -6 952 -4
rect 958 -6 960 -4
rect 972 -6 974 -4
rect 1004 -6 1006 -4
rect 1012 -6 1014 -4
rect 1027 -6 1029 -4
rect 1059 -6 1061 -4
rect 1067 -6 1069 -4
rect 1080 -6 1082 -4
rect 1112 -6 1114 -4
rect 1120 -6 1122 -4
<< pdifct0 >>
rect -273 329 -271 331
rect -263 350 -261 352
rect -263 343 -261 345
rect -247 336 -245 338
rect -247 329 -245 331
rect -227 344 -225 346
rect -202 350 -200 352
rect -190 331 -188 333
rect -167 350 -165 352
rect -167 343 -165 345
rect -155 342 -153 344
rect -155 335 -153 337
rect -145 350 -143 352
rect -145 343 -143 345
rect -113 350 -111 352
rect -113 343 -111 345
rect -103 342 -101 344
rect -103 335 -101 337
rect -91 350 -89 352
rect -91 343 -89 345
rect -56 350 -54 352
rect -68 331 -66 333
rect -34 343 -32 345
rect -15 350 -13 352
rect 9 343 11 345
rect 19 343 21 345
rect 19 336 21 338
rect 29 341 31 343
rect 49 343 51 345
rect 59 343 61 345
rect 59 336 61 338
rect 69 341 71 343
rect 100 350 102 352
rect 112 331 114 333
rect 135 350 137 352
rect 135 343 137 345
rect 147 342 149 344
rect 147 335 149 337
rect 157 350 159 352
rect 157 343 159 345
rect 189 350 191 352
rect 189 343 191 345
rect 199 342 201 344
rect 199 335 201 337
rect 211 350 213 352
rect 211 343 213 345
rect 246 350 248 352
rect 234 331 236 333
rect 268 343 270 345
rect 287 350 289 352
rect 316 343 318 345
rect 326 343 328 345
rect 326 336 328 338
rect 336 341 338 343
rect 377 350 379 352
rect 389 331 391 333
rect 412 350 414 352
rect 412 343 414 345
rect 424 342 426 344
rect 424 335 426 337
rect 434 350 436 352
rect 434 343 436 345
rect 466 350 468 352
rect 466 343 468 345
rect 476 342 478 344
rect 476 335 478 337
rect 488 350 490 352
rect 488 343 490 345
rect 523 350 525 352
rect 511 331 513 333
rect 545 343 547 345
rect 564 350 566 352
rect 593 343 595 345
rect 603 343 605 345
rect 603 336 605 338
rect 613 341 615 343
rect 653 350 655 352
rect 665 331 667 333
rect 688 350 690 352
rect 688 343 690 345
rect 700 342 702 344
rect 700 335 702 337
rect 710 350 712 352
rect 710 343 712 345
rect 742 350 744 352
rect 742 343 744 345
rect 752 342 754 344
rect 752 335 754 337
rect 764 350 766 352
rect 764 343 766 345
rect 799 350 801 352
rect 787 331 789 333
rect 821 343 823 345
rect 840 350 842 352
rect 869 343 871 345
rect 879 343 881 345
rect 879 336 881 338
rect 889 341 891 343
rect 930 350 932 352
rect 942 331 944 333
rect 965 350 967 352
rect 965 343 967 345
rect 977 342 979 344
rect 977 335 979 337
rect 987 350 989 352
rect 987 343 989 345
rect 1019 350 1021 352
rect 1019 343 1021 345
rect 1029 342 1031 344
rect 1029 335 1031 337
rect 1041 350 1043 352
rect 1041 343 1043 345
rect 1076 350 1078 352
rect 1064 331 1066 333
rect 1098 343 1100 345
rect 1117 350 1119 352
rect -273 245 -271 247
rect -263 231 -261 233
rect -247 245 -245 247
rect -247 238 -245 240
rect -263 224 -261 226
rect -227 230 -225 232
rect -190 243 -188 245
rect -202 224 -200 226
rect -167 231 -165 233
rect -167 224 -165 226
rect -155 239 -153 241
rect -155 232 -153 234
rect -145 231 -143 233
rect -145 224 -143 226
rect -113 231 -111 233
rect -113 224 -111 226
rect -103 239 -101 241
rect -103 232 -101 234
rect -91 231 -89 233
rect -91 224 -89 226
rect -68 243 -66 245
rect -56 224 -54 226
rect -34 231 -32 233
rect 9 231 11 233
rect 19 238 21 240
rect 19 231 21 233
rect 29 233 31 235
rect 49 231 51 233
rect -15 224 -13 226
rect 59 238 61 240
rect 59 231 61 233
rect 69 233 71 235
rect 112 243 114 245
rect 100 224 102 226
rect 135 231 137 233
rect 135 224 137 226
rect 147 239 149 241
rect 147 232 149 234
rect 157 231 159 233
rect 157 224 159 226
rect 189 231 191 233
rect 189 224 191 226
rect 199 239 201 241
rect 199 232 201 234
rect 211 231 213 233
rect 211 224 213 226
rect 234 243 236 245
rect 246 224 248 226
rect 268 231 270 233
rect 316 231 318 233
rect 326 238 328 240
rect 326 231 328 233
rect 336 233 338 235
rect 287 224 289 226
rect 389 243 391 245
rect 377 224 379 226
rect 412 231 414 233
rect 412 224 414 226
rect 424 239 426 241
rect 424 232 426 234
rect 434 231 436 233
rect 434 224 436 226
rect 466 231 468 233
rect 466 224 468 226
rect 476 239 478 241
rect 476 232 478 234
rect 488 231 490 233
rect 488 224 490 226
rect 511 243 513 245
rect 523 224 525 226
rect 545 231 547 233
rect 593 231 595 233
rect 603 238 605 240
rect 603 231 605 233
rect 613 233 615 235
rect 564 224 566 226
rect 665 243 667 245
rect 653 224 655 226
rect 688 231 690 233
rect 688 224 690 226
rect 700 239 702 241
rect 700 232 702 234
rect 710 231 712 233
rect 710 224 712 226
rect 742 231 744 233
rect 742 224 744 226
rect 752 239 754 241
rect 752 232 754 234
rect 764 231 766 233
rect 764 224 766 226
rect 787 243 789 245
rect 799 224 801 226
rect 821 231 823 233
rect 869 231 871 233
rect 879 238 881 240
rect 879 231 881 233
rect 889 233 891 235
rect 840 224 842 226
rect 942 243 944 245
rect 930 224 932 226
rect 965 231 967 233
rect 965 224 967 226
rect 977 239 979 241
rect 977 232 979 234
rect 987 231 989 233
rect 987 224 989 226
rect 1019 231 1021 233
rect 1019 224 1021 226
rect 1029 239 1031 241
rect 1029 232 1031 234
rect 1041 231 1043 233
rect 1041 224 1043 226
rect 1064 243 1066 245
rect 1076 224 1078 226
rect 1098 231 1100 233
rect 1117 224 1119 226
rect -273 185 -271 187
rect -263 206 -261 208
rect -263 199 -261 201
rect -247 192 -245 194
rect -247 185 -245 187
rect -227 200 -225 202
rect -202 206 -200 208
rect -190 187 -188 189
rect -167 206 -165 208
rect -167 199 -165 201
rect -155 198 -153 200
rect -155 191 -153 193
rect -145 206 -143 208
rect -145 199 -143 201
rect -113 206 -111 208
rect -113 199 -111 201
rect -103 198 -101 200
rect -103 191 -101 193
rect -91 206 -89 208
rect -91 199 -89 201
rect -56 206 -54 208
rect -68 187 -66 189
rect -34 199 -32 201
rect -15 206 -13 208
rect 9 199 11 201
rect 19 199 21 201
rect 19 192 21 194
rect 29 197 31 199
rect 49 199 51 201
rect 59 199 61 201
rect 59 192 61 194
rect 69 197 71 199
rect 100 206 102 208
rect 112 187 114 189
rect 135 206 137 208
rect 135 199 137 201
rect 147 198 149 200
rect 147 191 149 193
rect 157 206 159 208
rect 157 199 159 201
rect 189 206 191 208
rect 189 199 191 201
rect 199 198 201 200
rect 199 191 201 193
rect 211 206 213 208
rect 211 199 213 201
rect 246 206 248 208
rect 234 187 236 189
rect 268 199 270 201
rect 287 206 289 208
rect 316 199 318 201
rect 326 199 328 201
rect 326 192 328 194
rect 336 197 338 199
rect 377 206 379 208
rect 389 187 391 189
rect 412 206 414 208
rect 412 199 414 201
rect 424 198 426 200
rect 424 191 426 193
rect 434 206 436 208
rect 434 199 436 201
rect 466 206 468 208
rect 466 199 468 201
rect 476 198 478 200
rect 476 191 478 193
rect 488 206 490 208
rect 488 199 490 201
rect 523 206 525 208
rect 511 187 513 189
rect 545 199 547 201
rect 564 206 566 208
rect 593 199 595 201
rect 603 199 605 201
rect 603 192 605 194
rect 613 197 615 199
rect 653 206 655 208
rect 665 187 667 189
rect 688 206 690 208
rect 688 199 690 201
rect 700 198 702 200
rect 700 191 702 193
rect 710 206 712 208
rect 710 199 712 201
rect 742 206 744 208
rect 742 199 744 201
rect 752 198 754 200
rect 752 191 754 193
rect 764 206 766 208
rect 764 199 766 201
rect 799 206 801 208
rect 787 187 789 189
rect 821 199 823 201
rect 840 206 842 208
rect 869 199 871 201
rect 879 199 881 201
rect 879 192 881 194
rect 889 197 891 199
rect 930 206 932 208
rect 942 187 944 189
rect 965 206 967 208
rect 965 199 967 201
rect 977 198 979 200
rect 977 191 979 193
rect 987 206 989 208
rect 987 199 989 201
rect 1019 206 1021 208
rect 1019 199 1021 201
rect 1029 198 1031 200
rect 1029 191 1031 193
rect 1041 206 1043 208
rect 1041 199 1043 201
rect 1076 206 1078 208
rect 1064 187 1066 189
rect 1098 199 1100 201
rect 1117 206 1119 208
rect -273 101 -271 103
rect -263 87 -261 89
rect -247 101 -245 103
rect -247 94 -245 96
rect -263 80 -261 82
rect -227 86 -225 88
rect -190 99 -188 101
rect -202 80 -200 82
rect -167 87 -165 89
rect -167 80 -165 82
rect -155 95 -153 97
rect -155 88 -153 90
rect -145 87 -143 89
rect -145 80 -143 82
rect -113 87 -111 89
rect -113 80 -111 82
rect -103 95 -101 97
rect -103 88 -101 90
rect -91 87 -89 89
rect -91 80 -89 82
rect -68 99 -66 101
rect -56 80 -54 82
rect -34 87 -32 89
rect 9 87 11 89
rect 19 94 21 96
rect 19 87 21 89
rect 29 89 31 91
rect 49 87 51 89
rect -15 80 -13 82
rect 59 94 61 96
rect 59 87 61 89
rect 69 89 71 91
rect 112 99 114 101
rect 100 80 102 82
rect 135 87 137 89
rect 135 80 137 82
rect 147 95 149 97
rect 147 88 149 90
rect 157 87 159 89
rect 157 80 159 82
rect 189 87 191 89
rect 189 80 191 82
rect 199 95 201 97
rect 199 88 201 90
rect 211 87 213 89
rect 211 80 213 82
rect 234 99 236 101
rect 246 80 248 82
rect 268 87 270 89
rect 316 87 318 89
rect 326 94 328 96
rect 326 87 328 89
rect 336 89 338 91
rect 287 80 289 82
rect 389 99 391 101
rect 377 80 379 82
rect 412 87 414 89
rect 412 80 414 82
rect 424 95 426 97
rect 424 88 426 90
rect 434 87 436 89
rect 434 80 436 82
rect 466 87 468 89
rect 466 80 468 82
rect 476 95 478 97
rect 476 88 478 90
rect 488 87 490 89
rect 488 80 490 82
rect 511 99 513 101
rect 523 80 525 82
rect 545 87 547 89
rect 593 87 595 89
rect 603 94 605 96
rect 603 87 605 89
rect 613 89 615 91
rect 564 80 566 82
rect 665 99 667 101
rect 653 80 655 82
rect 688 87 690 89
rect 688 80 690 82
rect 700 95 702 97
rect 700 88 702 90
rect 710 87 712 89
rect 710 80 712 82
rect 742 87 744 89
rect 742 80 744 82
rect 752 95 754 97
rect 752 88 754 90
rect 764 87 766 89
rect 764 80 766 82
rect 787 99 789 101
rect 799 80 801 82
rect 821 87 823 89
rect 869 87 871 89
rect 879 94 881 96
rect 879 87 881 89
rect 889 89 891 91
rect 840 80 842 82
rect 942 99 944 101
rect 930 80 932 82
rect 965 87 967 89
rect 965 80 967 82
rect 977 95 979 97
rect 977 88 979 90
rect 987 87 989 89
rect 987 80 989 82
rect 1019 87 1021 89
rect 1019 80 1021 82
rect 1029 95 1031 97
rect 1029 88 1031 90
rect 1041 87 1043 89
rect 1041 80 1043 82
rect 1064 99 1066 101
rect 1076 80 1078 82
rect 1098 87 1100 89
rect 1117 80 1119 82
rect -273 41 -271 43
rect -263 62 -261 64
rect -263 55 -261 57
rect -247 48 -245 50
rect -247 41 -245 43
rect -227 56 -225 58
rect -202 62 -200 64
rect -190 43 -188 45
rect -167 62 -165 64
rect -167 55 -165 57
rect -155 54 -153 56
rect -155 47 -153 49
rect -145 62 -143 64
rect -145 55 -143 57
rect -113 62 -111 64
rect -113 55 -111 57
rect -103 54 -101 56
rect -103 47 -101 49
rect -91 62 -89 64
rect -91 55 -89 57
rect -56 62 -54 64
rect -68 43 -66 45
rect -34 55 -32 57
rect -15 62 -13 64
rect 9 55 11 57
rect 19 55 21 57
rect 19 48 21 50
rect 29 53 31 55
rect 49 55 51 57
rect 59 55 61 57
rect 59 48 61 50
rect 69 53 71 55
rect 100 62 102 64
rect 112 43 114 45
rect 135 62 137 64
rect 135 55 137 57
rect 147 54 149 56
rect 147 47 149 49
rect 157 62 159 64
rect 157 55 159 57
rect 189 62 191 64
rect 189 55 191 57
rect 199 54 201 56
rect 199 47 201 49
rect 211 62 213 64
rect 211 55 213 57
rect 246 62 248 64
rect 234 43 236 45
rect 268 55 270 57
rect 287 62 289 64
rect 316 55 318 57
rect 326 55 328 57
rect 326 48 328 50
rect 336 53 338 55
rect 377 62 379 64
rect 389 43 391 45
rect 412 62 414 64
rect 412 55 414 57
rect 424 54 426 56
rect 424 47 426 49
rect 434 62 436 64
rect 434 55 436 57
rect 466 62 468 64
rect 466 55 468 57
rect 476 54 478 56
rect 476 47 478 49
rect 488 62 490 64
rect 488 55 490 57
rect 523 62 525 64
rect 511 43 513 45
rect 545 55 547 57
rect 564 62 566 64
rect 593 55 595 57
rect 603 55 605 57
rect 603 48 605 50
rect 613 53 615 55
rect 653 62 655 64
rect 665 43 667 45
rect 688 62 690 64
rect 688 55 690 57
rect 700 54 702 56
rect 700 47 702 49
rect 710 62 712 64
rect 710 55 712 57
rect 742 62 744 64
rect 742 55 744 57
rect 752 54 754 56
rect 752 47 754 49
rect 764 62 766 64
rect 764 55 766 57
rect 799 62 801 64
rect 787 43 789 45
rect 821 55 823 57
rect 840 62 842 64
rect 869 55 871 57
rect 879 55 881 57
rect 879 48 881 50
rect 889 53 891 55
rect 930 62 932 64
rect 942 43 944 45
rect 965 62 967 64
rect 965 55 967 57
rect 977 54 979 56
rect 977 47 979 49
rect 987 62 989 64
rect 987 55 989 57
rect 1019 62 1021 64
rect 1019 55 1021 57
rect 1029 54 1031 56
rect 1029 47 1031 49
rect 1041 62 1043 64
rect 1041 55 1043 57
rect 1076 62 1078 64
rect 1064 43 1066 45
rect 1098 55 1100 57
rect 1117 62 1119 64
rect -134 -49 -132 -47
rect -112 -55 -110 -53
rect -82 -49 -80 -47
rect -60 -55 -58 -53
rect -30 -49 -28 -47
rect -8 -55 -6 -53
rect 22 -49 24 -47
rect 44 -55 46 -53
rect 74 -49 76 -47
rect 96 -55 98 -53
rect 127 -49 129 -47
rect 149 -55 151 -53
rect 315 -49 317 -47
rect 337 -55 339 -53
rect 368 -49 370 -47
rect 390 -55 392 -53
rect 420 -49 422 -47
rect 442 -55 444 -53
rect 472 -49 474 -47
rect 494 -55 496 -53
rect 524 -49 526 -47
rect 546 -55 548 -53
rect 623 -49 625 -47
rect 645 -55 647 -53
rect 676 -49 678 -47
rect 698 -55 700 -53
rect 728 -49 730 -47
rect 750 -55 752 -53
rect 780 -49 782 -47
rect 802 -55 804 -53
rect 832 -49 834 -47
rect 854 -55 856 -53
rect 884 -49 886 -47
rect 906 -55 908 -53
rect 937 -49 939 -47
rect 959 -55 961 -53
rect 991 -49 993 -47
rect 1013 -55 1015 -53
rect 1046 -49 1048 -47
rect 1068 -55 1070 -53
rect 1099 -49 1101 -47
rect 1121 -55 1123 -53
<< pdifct1 >>
rect -237 336 -235 338
rect -213 338 -211 340
rect -213 331 -211 333
rect -135 335 -133 337
rect -135 328 -133 330
rect -123 335 -121 337
rect -123 328 -121 330
rect -45 338 -43 340
rect -45 331 -43 333
rect -4 340 -2 342
rect -4 333 -2 335
rect 39 336 41 338
rect 39 329 41 331
rect 79 336 81 338
rect 79 329 81 331
rect 89 338 91 340
rect 89 331 91 333
rect 167 335 169 337
rect 167 328 169 330
rect 179 335 181 337
rect 179 328 181 330
rect 257 338 259 340
rect 257 331 259 333
rect 298 340 300 342
rect 298 333 300 335
rect 346 336 348 338
rect 346 329 348 331
rect 366 338 368 340
rect 366 331 368 333
rect 444 335 446 337
rect 444 328 446 330
rect 456 335 458 337
rect 456 328 458 330
rect 534 338 536 340
rect 534 331 536 333
rect 575 340 577 342
rect 575 333 577 335
rect 623 336 625 338
rect 623 329 625 331
rect 642 338 644 340
rect 642 331 644 333
rect 720 335 722 337
rect 720 328 722 330
rect 732 335 734 337
rect 732 328 734 330
rect 810 338 812 340
rect 810 331 812 333
rect 851 340 853 342
rect 851 333 853 335
rect 899 336 901 338
rect 899 329 901 331
rect 919 338 921 340
rect 919 331 921 333
rect 997 335 999 337
rect 997 328 999 330
rect 1009 335 1011 337
rect 1009 328 1011 330
rect 1087 338 1089 340
rect 1087 331 1089 333
rect 1128 340 1130 342
rect 1128 333 1130 335
rect -237 238 -235 240
rect -213 243 -211 245
rect -213 236 -211 238
rect -135 246 -133 248
rect -135 239 -133 241
rect -123 246 -121 248
rect -123 239 -121 241
rect -45 243 -43 245
rect -45 236 -43 238
rect -4 241 -2 243
rect -4 234 -2 236
rect 39 244 41 246
rect 39 236 41 238
rect 79 245 81 247
rect 79 238 81 240
rect 89 243 91 245
rect 89 236 91 238
rect 167 246 169 248
rect 167 239 169 241
rect 179 246 181 248
rect 179 239 181 241
rect 257 243 259 245
rect 257 236 259 238
rect 298 241 300 243
rect 298 234 300 236
rect 346 245 348 247
rect 346 238 348 240
rect 366 243 368 245
rect 366 236 368 238
rect 444 246 446 248
rect 444 239 446 241
rect 456 246 458 248
rect 456 239 458 241
rect 534 243 536 245
rect 534 236 536 238
rect 575 241 577 243
rect 575 234 577 236
rect 623 245 625 247
rect 623 238 625 240
rect 642 243 644 245
rect 642 236 644 238
rect 720 246 722 248
rect 720 239 722 241
rect 732 246 734 248
rect 732 239 734 241
rect 810 243 812 245
rect 810 236 812 238
rect 851 241 853 243
rect 851 234 853 236
rect 899 245 901 247
rect 899 238 901 240
rect 919 243 921 245
rect 919 236 921 238
rect 997 246 999 248
rect 997 239 999 241
rect 1009 246 1011 248
rect 1009 239 1011 241
rect 1087 243 1089 245
rect 1087 236 1089 238
rect 1128 241 1130 243
rect 1128 234 1130 236
rect -237 192 -235 194
rect -213 194 -211 196
rect -213 187 -211 189
rect -135 191 -133 193
rect -135 184 -133 186
rect -123 191 -121 193
rect -123 184 -121 186
rect -45 194 -43 196
rect -45 187 -43 189
rect -4 196 -2 198
rect -4 189 -2 191
rect 39 195 41 197
rect 39 187 41 189
rect 79 192 81 194
rect 79 185 81 187
rect 89 194 91 196
rect 89 187 91 189
rect 167 191 169 193
rect 167 184 169 186
rect 179 191 181 193
rect 179 184 181 186
rect 257 194 259 196
rect 257 187 259 189
rect 298 196 300 198
rect 298 189 300 191
rect 346 192 348 194
rect 346 185 348 187
rect 366 194 368 196
rect 366 187 368 189
rect 444 191 446 193
rect 444 184 446 186
rect 456 191 458 193
rect 456 184 458 186
rect 534 194 536 196
rect 534 187 536 189
rect 575 196 577 198
rect 575 189 577 191
rect 623 192 625 194
rect 623 185 625 187
rect 642 194 644 196
rect 642 187 644 189
rect 720 191 722 193
rect 720 184 722 186
rect 732 191 734 193
rect 732 184 734 186
rect 810 194 812 196
rect 810 187 812 189
rect 851 196 853 198
rect 851 189 853 191
rect 899 192 901 194
rect 899 185 901 187
rect 919 194 921 196
rect 919 187 921 189
rect 997 191 999 193
rect 997 184 999 186
rect 1009 191 1011 193
rect 1009 184 1011 186
rect 1087 194 1089 196
rect 1087 187 1089 189
rect 1128 196 1130 198
rect 1128 189 1130 191
rect -237 94 -235 96
rect -213 99 -211 101
rect -213 92 -211 94
rect -135 102 -133 104
rect -135 95 -133 97
rect -123 102 -121 104
rect -123 95 -121 97
rect -45 99 -43 101
rect -45 92 -43 94
rect -4 97 -2 99
rect -4 90 -2 92
rect 39 98 41 100
rect 39 91 41 93
rect 79 101 81 103
rect 79 94 81 96
rect 89 99 91 101
rect 89 92 91 94
rect 167 102 169 104
rect 167 95 169 97
rect 179 102 181 104
rect 179 95 181 97
rect 257 99 259 101
rect 257 92 259 94
rect 298 97 300 99
rect 298 90 300 92
rect 346 101 348 103
rect 346 94 348 96
rect 366 99 368 101
rect 366 92 368 94
rect 444 102 446 104
rect 444 95 446 97
rect 456 102 458 104
rect 456 95 458 97
rect 534 99 536 101
rect 534 92 536 94
rect 575 97 577 99
rect 575 90 577 92
rect 623 101 625 103
rect 623 94 625 96
rect 642 99 644 101
rect 642 92 644 94
rect 720 102 722 104
rect 720 95 722 97
rect 732 102 734 104
rect 732 95 734 97
rect 810 99 812 101
rect 810 92 812 94
rect 851 97 853 99
rect 851 90 853 92
rect 899 101 901 103
rect 899 94 901 96
rect 919 99 921 101
rect 919 92 921 94
rect 997 102 999 104
rect 997 95 999 97
rect 1009 102 1011 104
rect 1009 95 1011 97
rect 1087 99 1089 101
rect 1087 92 1089 94
rect 1128 97 1130 99
rect 1128 90 1130 92
rect -237 48 -235 50
rect -213 50 -211 52
rect -213 43 -211 45
rect -135 47 -133 49
rect -135 40 -133 42
rect -123 47 -121 49
rect -123 40 -121 42
rect -45 50 -43 52
rect -45 43 -43 45
rect -4 52 -2 54
rect -4 45 -2 47
rect 39 48 41 50
rect 39 41 41 43
rect 79 48 81 50
rect 79 41 81 43
rect 89 50 91 52
rect 89 43 91 45
rect 167 47 169 49
rect 167 40 169 42
rect 179 47 181 49
rect 179 40 181 42
rect 257 50 259 52
rect 257 43 259 45
rect 298 52 300 54
rect 298 45 300 47
rect 346 48 348 50
rect 346 41 348 43
rect 366 50 368 52
rect 366 43 368 45
rect 444 47 446 49
rect 444 40 446 42
rect 456 47 458 49
rect 456 40 458 42
rect 534 50 536 52
rect 534 43 536 45
rect 575 52 577 54
rect 575 45 577 47
rect 623 48 625 50
rect 623 41 625 43
rect 642 50 644 52
rect 642 43 644 45
rect 720 47 722 49
rect 720 40 722 42
rect 732 47 734 49
rect 732 40 734 42
rect 810 50 812 52
rect 810 43 812 45
rect 851 52 853 54
rect 851 45 853 47
rect 899 48 901 50
rect 899 41 901 43
rect 919 50 921 52
rect 919 43 921 45
rect 997 47 999 49
rect 997 40 999 42
rect 1009 47 1011 49
rect 1009 40 1011 42
rect 1087 50 1089 52
rect 1087 43 1089 45
rect 1128 52 1130 54
rect 1128 45 1130 47
rect -154 -55 -152 -53
rect -102 -55 -100 -53
rect -143 -66 -141 -64
rect -50 -55 -48 -53
rect -123 -66 -121 -64
rect -91 -66 -89 -64
rect 2 -55 4 -53
rect -71 -66 -69 -64
rect -39 -66 -37 -64
rect 54 -55 56 -53
rect -19 -66 -17 -64
rect 13 -66 15 -64
rect 107 -55 109 -53
rect 33 -66 35 -64
rect 65 -66 67 -64
rect 174 -41 176 -39
rect 194 -41 196 -39
rect 214 -41 216 -39
rect 236 -41 238 -39
rect 258 -41 260 -39
rect 280 -41 282 -39
rect 85 -66 87 -64
rect 118 -66 120 -64
rect 295 -55 297 -53
rect 138 -66 140 -64
rect 164 -66 166 -64
rect 184 -66 186 -64
rect 204 -66 206 -64
rect 226 -66 228 -64
rect 248 -66 250 -64
rect 270 -66 272 -64
rect 348 -55 350 -53
rect 306 -66 308 -64
rect 400 -55 402 -53
rect 326 -66 328 -64
rect 359 -66 361 -64
rect 452 -55 454 -53
rect 379 -66 381 -64
rect 411 -66 413 -64
rect 504 -55 506 -53
rect 431 -66 433 -64
rect 463 -66 465 -64
rect 569 -41 571 -39
rect 590 -41 592 -39
rect 483 -66 485 -64
rect 515 -66 517 -64
rect 603 -55 605 -53
rect 535 -66 537 -64
rect 559 -66 561 -64
rect 580 -66 582 -64
rect 656 -55 658 -53
rect 614 -66 616 -64
rect 708 -55 710 -53
rect 634 -66 636 -64
rect 667 -66 669 -64
rect 760 -55 762 -53
rect 687 -66 689 -64
rect 719 -66 721 -64
rect 812 -55 814 -53
rect 739 -66 741 -64
rect 771 -66 773 -64
rect 864 -55 866 -53
rect 791 -66 793 -64
rect 823 -66 825 -64
rect 917 -55 919 -53
rect 843 -66 845 -64
rect 875 -66 877 -64
rect 971 -55 973 -53
rect 895 -66 897 -64
rect 928 -66 930 -64
rect 1026 -55 1028 -53
rect 948 -66 950 -64
rect 982 -66 984 -64
rect 1079 -55 1081 -53
rect 1002 -66 1004 -64
rect 1037 -66 1039 -64
rect 1057 -66 1059 -64
rect 1090 -66 1092 -64
rect 1110 -66 1112 -64
<< alu0 >>
rect -264 350 -263 352
rect -261 350 -260 352
rect -264 345 -260 350
rect -204 350 -202 352
rect -200 350 -198 352
rect -204 349 -198 350
rect -169 350 -167 352
rect -165 350 -163 352
rect -264 343 -263 345
rect -261 343 -260 345
rect -264 341 -260 343
rect -256 346 -223 347
rect -256 344 -227 346
rect -225 344 -223 346
rect -256 343 -223 344
rect -169 345 -163 350
rect -147 350 -145 352
rect -143 350 -141 352
rect -169 343 -167 345
rect -165 343 -163 345
rect -256 332 -252 343
rect -169 342 -163 343
rect -156 344 -152 346
rect -156 342 -155 344
rect -153 342 -152 344
rect -147 345 -141 350
rect -147 343 -145 345
rect -143 343 -141 345
rect -147 342 -141 343
rect -115 350 -113 352
rect -111 350 -109 352
rect -115 345 -109 350
rect -93 350 -91 352
rect -89 350 -87 352
rect -115 343 -113 345
rect -111 343 -109 345
rect -115 342 -109 343
rect -104 344 -100 346
rect -104 342 -103 344
rect -101 342 -100 344
rect -93 345 -87 350
rect -58 350 -56 352
rect -54 350 -52 352
rect -58 349 -52 350
rect -17 350 -15 352
rect -13 350 -11 352
rect -17 349 -11 350
rect -93 343 -91 345
rect -89 343 -87 345
rect -93 342 -87 343
rect -36 345 -19 346
rect -36 343 -34 345
rect -32 343 -19 345
rect -36 342 -19 343
rect 7 345 13 352
rect 7 343 9 345
rect 11 343 13 345
rect 7 342 13 343
rect 18 345 22 347
rect 18 343 19 345
rect 21 343 22 345
rect -275 331 -252 332
rect -275 329 -273 331
rect -271 329 -252 331
rect -275 328 -252 329
rect -275 322 -271 328
rect -282 318 -271 322
rect -282 312 -278 318
rect -256 322 -252 328
rect -248 338 -244 340
rect -248 336 -247 338
rect -245 336 -244 338
rect -248 331 -244 336
rect -248 329 -247 331
rect -245 330 -244 331
rect -245 329 -232 330
rect -248 326 -232 329
rect -236 324 -232 326
rect -236 322 -231 324
rect -256 321 -240 322
rect -256 319 -244 321
rect -242 319 -240 321
rect -256 318 -240 319
rect -236 320 -234 322
rect -232 320 -231 322
rect -236 318 -231 320
rect -282 310 -281 312
rect -279 310 -278 312
rect -282 308 -278 310
rect -236 314 -232 318
rect -256 310 -232 314
rect -256 307 -252 310
rect -256 305 -255 307
rect -253 305 -252 307
rect -269 304 -263 305
rect -269 302 -267 304
rect -265 302 -263 304
rect -256 303 -252 305
rect -199 338 -175 342
rect -156 338 -152 342
rect -201 334 -195 338
rect -179 337 -139 338
rect -179 335 -155 337
rect -153 335 -139 337
rect -201 324 -197 334
rect -191 333 -187 335
rect -179 334 -139 335
rect -191 331 -190 333
rect -188 331 -187 333
rect -191 330 -187 331
rect -201 322 -200 324
rect -198 322 -197 324
rect -201 320 -197 322
rect -194 326 -187 330
rect -194 315 -190 326
rect -151 321 -147 326
rect -151 319 -150 321
rect -148 319 -147 321
rect -208 314 -190 315
rect -208 312 -206 314
rect -204 313 -190 314
rect -204 312 -179 313
rect -208 311 -183 312
rect -194 310 -183 311
rect -181 310 -179 312
rect -194 309 -179 310
rect -174 312 -170 314
rect -174 310 -173 312
rect -171 310 -170 312
rect -174 305 -170 310
rect -151 317 -147 319
rect -143 323 -139 334
rect -143 321 -137 323
rect -143 319 -140 321
rect -138 319 -137 321
rect -143 317 -137 319
rect -143 314 -139 317
rect -159 310 -139 314
rect -159 306 -155 310
rect -195 304 -173 305
rect -269 296 -263 302
rect -204 301 -200 303
rect -195 302 -193 304
rect -191 303 -173 304
rect -171 303 -170 305
rect -191 302 -170 303
rect -165 305 -155 306
rect -165 303 -163 305
rect -161 303 -155 305
rect -165 302 -155 303
rect -104 338 -100 342
rect -81 338 -57 342
rect -117 337 -77 338
rect -117 335 -103 337
rect -101 335 -77 337
rect -117 334 -77 335
rect -117 323 -113 334
rect -69 333 -65 335
rect -61 334 -55 338
rect -69 331 -68 333
rect -66 331 -65 333
rect -69 330 -65 331
rect -69 326 -62 330
rect -119 321 -113 323
rect -119 319 -118 321
rect -116 319 -113 321
rect -119 317 -113 319
rect -109 321 -105 326
rect -109 319 -108 321
rect -106 319 -105 321
rect -109 317 -105 319
rect -117 314 -113 317
rect -117 310 -97 314
rect -101 306 -97 310
rect -66 315 -62 326
rect -59 324 -55 334
rect -59 322 -58 324
rect -56 322 -55 324
rect -59 320 -55 322
rect -66 314 -48 315
rect -86 312 -82 314
rect -66 313 -52 314
rect -86 310 -85 312
rect -83 310 -82 312
rect -101 305 -91 306
rect -101 303 -95 305
rect -93 303 -91 305
rect -101 302 -91 303
rect -86 305 -82 310
rect -77 312 -52 313
rect -50 312 -48 314
rect -77 310 -75 312
rect -73 311 -48 312
rect -73 310 -62 311
rect -77 309 -62 310
rect -23 338 -19 342
rect -23 334 -8 338
rect -33 325 -27 326
rect -12 321 -8 334
rect -5 331 -4 342
rect -12 319 -11 321
rect -9 319 -8 321
rect -12 313 -8 319
rect 18 338 22 343
rect 27 343 33 352
rect 27 341 29 343
rect 31 341 33 343
rect 47 345 53 352
rect 47 343 49 345
rect 51 343 53 345
rect 47 342 53 343
rect 58 345 62 347
rect 58 343 59 345
rect 61 343 62 345
rect 27 340 33 341
rect 18 336 19 338
rect 21 337 22 338
rect 21 336 35 337
rect 18 333 35 336
rect -26 312 -8 313
rect -26 310 -24 312
rect -22 310 -8 312
rect -26 309 -8 310
rect 31 321 35 333
rect 31 319 32 321
rect 34 319 35 321
rect 31 314 35 319
rect 23 310 35 314
rect 58 338 62 343
rect 67 343 73 352
rect 98 350 100 352
rect 102 350 104 352
rect 98 349 104 350
rect 133 350 135 352
rect 137 350 139 352
rect 67 341 69 343
rect 71 341 73 343
rect 133 345 139 350
rect 155 350 157 352
rect 159 350 161 352
rect 133 343 135 345
rect 137 343 139 345
rect 133 342 139 343
rect 146 344 150 346
rect 146 342 147 344
rect 149 342 150 344
rect 155 345 161 350
rect 155 343 157 345
rect 159 343 161 345
rect 155 342 161 343
rect 187 350 189 352
rect 191 350 193 352
rect 187 345 193 350
rect 209 350 211 352
rect 213 350 215 352
rect 187 343 189 345
rect 191 343 193 345
rect 187 342 193 343
rect 198 344 202 346
rect 198 342 199 344
rect 201 342 202 344
rect 209 345 215 350
rect 244 350 246 352
rect 248 350 250 352
rect 244 349 250 350
rect 285 350 287 352
rect 289 350 291 352
rect 285 349 291 350
rect 209 343 211 345
rect 213 343 215 345
rect 209 342 215 343
rect 266 345 283 346
rect 266 343 268 345
rect 270 343 283 345
rect 266 342 283 343
rect 314 345 320 352
rect 314 343 316 345
rect 318 343 320 345
rect 314 342 320 343
rect 325 345 329 347
rect 325 343 326 345
rect 328 343 329 345
rect 67 340 73 341
rect 58 336 59 338
rect 61 337 62 338
rect 61 336 75 337
rect 58 333 75 336
rect 23 306 27 310
rect 38 307 39 309
rect 71 321 75 333
rect 71 319 72 321
rect 74 319 75 321
rect 71 314 75 319
rect 63 310 75 314
rect -86 303 -85 305
rect -83 304 -61 305
rect -83 303 -65 304
rect -86 302 -65 303
rect -63 302 -61 304
rect -195 301 -170 302
rect -86 301 -61 302
rect -56 301 -52 303
rect 7 305 27 306
rect 7 303 9 305
rect 11 303 27 305
rect 7 302 27 303
rect 63 306 67 310
rect 78 307 79 309
rect 47 305 67 306
rect 47 303 49 305
rect 51 303 67 305
rect 47 302 67 303
rect 103 338 127 342
rect 146 338 150 342
rect 101 334 107 338
rect 123 337 163 338
rect 123 335 147 337
rect 149 335 163 337
rect 101 324 105 334
rect 111 333 115 335
rect 123 334 163 335
rect 111 331 112 333
rect 114 331 115 333
rect 111 330 115 331
rect 101 322 102 324
rect 104 322 105 324
rect 101 320 105 322
rect 108 326 115 330
rect 108 315 112 326
rect 151 321 155 326
rect 151 319 152 321
rect 154 319 155 321
rect 94 314 112 315
rect 94 312 96 314
rect 98 313 112 314
rect 98 312 123 313
rect 94 311 119 312
rect 108 310 119 311
rect 121 310 123 312
rect 108 309 123 310
rect 128 312 132 314
rect 128 310 129 312
rect 131 310 132 312
rect 128 305 132 310
rect 151 317 155 319
rect 159 323 163 334
rect 159 321 165 323
rect 159 319 162 321
rect 164 319 165 321
rect 159 317 165 319
rect 159 314 163 317
rect 143 310 163 314
rect 143 306 147 310
rect 107 304 129 305
rect 98 301 102 303
rect 107 302 109 304
rect 111 303 129 304
rect 131 303 132 305
rect 111 302 132 303
rect 137 305 147 306
rect 137 303 139 305
rect 141 303 147 305
rect 137 302 147 303
rect 198 338 202 342
rect 221 338 245 342
rect 185 337 225 338
rect 185 335 199 337
rect 201 335 225 337
rect 185 334 225 335
rect 185 323 189 334
rect 233 333 237 335
rect 241 334 247 338
rect 233 331 234 333
rect 236 331 237 333
rect 233 330 237 331
rect 233 326 240 330
rect 183 321 189 323
rect 183 319 184 321
rect 186 319 189 321
rect 183 317 189 319
rect 193 321 197 326
rect 193 319 194 321
rect 196 319 197 321
rect 193 317 197 319
rect 185 314 189 317
rect 185 310 205 314
rect 201 306 205 310
rect 236 315 240 326
rect 243 324 247 334
rect 243 322 244 324
rect 246 322 247 324
rect 243 320 247 322
rect 236 314 254 315
rect 216 312 220 314
rect 236 313 250 314
rect 216 310 217 312
rect 219 310 220 312
rect 201 305 211 306
rect 201 303 207 305
rect 209 303 211 305
rect 201 302 211 303
rect 216 305 220 310
rect 225 312 250 313
rect 252 312 254 314
rect 225 310 227 312
rect 229 311 254 312
rect 229 310 240 311
rect 225 309 240 310
rect 279 338 283 342
rect 279 334 294 338
rect 269 325 275 326
rect 290 321 294 334
rect 297 331 298 342
rect 290 319 291 321
rect 293 319 294 321
rect 290 313 294 319
rect 325 338 329 343
rect 334 343 340 352
rect 375 350 377 352
rect 379 350 381 352
rect 375 349 381 350
rect 410 350 412 352
rect 414 350 416 352
rect 334 341 336 343
rect 338 341 340 343
rect 410 345 416 350
rect 432 350 434 352
rect 436 350 438 352
rect 410 343 412 345
rect 414 343 416 345
rect 410 342 416 343
rect 423 344 427 346
rect 423 342 424 344
rect 426 342 427 344
rect 432 345 438 350
rect 432 343 434 345
rect 436 343 438 345
rect 432 342 438 343
rect 464 350 466 352
rect 468 350 470 352
rect 464 345 470 350
rect 486 350 488 352
rect 490 350 492 352
rect 464 343 466 345
rect 468 343 470 345
rect 464 342 470 343
rect 475 344 479 346
rect 475 342 476 344
rect 478 342 479 344
rect 486 345 492 350
rect 521 350 523 352
rect 525 350 527 352
rect 521 349 527 350
rect 562 350 564 352
rect 566 350 568 352
rect 562 349 568 350
rect 486 343 488 345
rect 490 343 492 345
rect 486 342 492 343
rect 543 345 560 346
rect 543 343 545 345
rect 547 343 560 345
rect 543 342 560 343
rect 591 345 597 352
rect 591 343 593 345
rect 595 343 597 345
rect 591 342 597 343
rect 602 345 606 347
rect 602 343 603 345
rect 605 343 606 345
rect 334 340 340 341
rect 325 336 326 338
rect 328 337 329 338
rect 328 336 342 337
rect 325 333 342 336
rect 276 312 294 313
rect 276 310 278 312
rect 280 310 294 312
rect 276 309 294 310
rect 338 321 342 333
rect 338 319 339 321
rect 341 319 342 321
rect 338 314 342 319
rect 330 310 342 314
rect 330 306 334 310
rect 345 307 346 309
rect 216 303 217 305
rect 219 304 241 305
rect 219 303 237 304
rect 216 302 237 303
rect 239 302 241 304
rect 107 301 132 302
rect 216 301 241 302
rect 246 301 250 303
rect 314 305 334 306
rect 314 303 316 305
rect 318 303 334 305
rect 314 302 334 303
rect 380 338 404 342
rect 423 338 427 342
rect 378 334 384 338
rect 400 337 440 338
rect 400 335 424 337
rect 426 335 440 337
rect 378 324 382 334
rect 388 333 392 335
rect 400 334 440 335
rect 388 331 389 333
rect 391 331 392 333
rect 388 330 392 331
rect 378 322 379 324
rect 381 322 382 324
rect 378 320 382 322
rect 385 326 392 330
rect 385 315 389 326
rect 428 321 432 326
rect 428 319 429 321
rect 431 319 432 321
rect 371 314 389 315
rect 371 312 373 314
rect 375 313 389 314
rect 375 312 400 313
rect 371 311 396 312
rect 385 310 396 311
rect 398 310 400 312
rect 385 309 400 310
rect 405 312 409 314
rect 405 310 406 312
rect 408 310 409 312
rect 405 305 409 310
rect 428 317 432 319
rect 436 323 440 334
rect 436 321 442 323
rect 436 319 439 321
rect 441 319 442 321
rect 436 317 442 319
rect 436 314 440 317
rect 420 310 440 314
rect 420 306 424 310
rect 384 304 406 305
rect 375 301 379 303
rect 384 302 386 304
rect 388 303 406 304
rect 408 303 409 305
rect 388 302 409 303
rect 414 305 424 306
rect 414 303 416 305
rect 418 303 424 305
rect 414 302 424 303
rect 475 338 479 342
rect 498 338 522 342
rect 462 337 502 338
rect 462 335 476 337
rect 478 335 502 337
rect 462 334 502 335
rect 462 323 466 334
rect 510 333 514 335
rect 518 334 524 338
rect 510 331 511 333
rect 513 331 514 333
rect 510 330 514 331
rect 510 326 517 330
rect 460 321 466 323
rect 460 319 461 321
rect 463 319 466 321
rect 460 317 466 319
rect 470 321 474 326
rect 470 319 471 321
rect 473 319 474 321
rect 470 317 474 319
rect 462 314 466 317
rect 462 310 482 314
rect 478 306 482 310
rect 513 315 517 326
rect 520 324 524 334
rect 520 322 521 324
rect 523 322 524 324
rect 520 320 524 322
rect 513 314 531 315
rect 493 312 497 314
rect 513 313 527 314
rect 493 310 494 312
rect 496 310 497 312
rect 478 305 488 306
rect 478 303 484 305
rect 486 303 488 305
rect 478 302 488 303
rect 493 305 497 310
rect 502 312 527 313
rect 529 312 531 314
rect 502 310 504 312
rect 506 311 531 312
rect 506 310 517 311
rect 502 309 517 310
rect 556 338 560 342
rect 556 334 571 338
rect 546 325 552 326
rect 567 321 571 334
rect 574 331 575 342
rect 567 319 568 321
rect 570 319 571 321
rect 567 313 571 319
rect 602 338 606 343
rect 611 343 617 352
rect 651 350 653 352
rect 655 350 657 352
rect 651 349 657 350
rect 686 350 688 352
rect 690 350 692 352
rect 611 341 613 343
rect 615 341 617 343
rect 686 345 692 350
rect 708 350 710 352
rect 712 350 714 352
rect 686 343 688 345
rect 690 343 692 345
rect 686 342 692 343
rect 699 344 703 346
rect 699 342 700 344
rect 702 342 703 344
rect 708 345 714 350
rect 708 343 710 345
rect 712 343 714 345
rect 708 342 714 343
rect 740 350 742 352
rect 744 350 746 352
rect 740 345 746 350
rect 762 350 764 352
rect 766 350 768 352
rect 740 343 742 345
rect 744 343 746 345
rect 740 342 746 343
rect 751 344 755 346
rect 751 342 752 344
rect 754 342 755 344
rect 762 345 768 350
rect 797 350 799 352
rect 801 350 803 352
rect 797 349 803 350
rect 838 350 840 352
rect 842 350 844 352
rect 838 349 844 350
rect 762 343 764 345
rect 766 343 768 345
rect 762 342 768 343
rect 819 345 836 346
rect 819 343 821 345
rect 823 343 836 345
rect 819 342 836 343
rect 867 345 873 352
rect 867 343 869 345
rect 871 343 873 345
rect 867 342 873 343
rect 878 345 882 347
rect 878 343 879 345
rect 881 343 882 345
rect 611 340 617 341
rect 602 336 603 338
rect 605 337 606 338
rect 605 336 619 337
rect 602 333 619 336
rect 553 312 571 313
rect 553 310 555 312
rect 557 310 571 312
rect 553 309 571 310
rect 615 321 619 333
rect 615 319 616 321
rect 618 319 619 321
rect 615 314 619 319
rect 607 310 619 314
rect 607 306 611 310
rect 622 307 623 309
rect 493 303 494 305
rect 496 304 518 305
rect 496 303 514 304
rect 493 302 514 303
rect 516 302 518 304
rect 384 301 409 302
rect 493 301 518 302
rect 523 301 527 303
rect 591 305 611 306
rect 591 303 593 305
rect 595 303 611 305
rect 591 302 611 303
rect 656 338 680 342
rect 699 338 703 342
rect 654 334 660 338
rect 676 337 716 338
rect 676 335 700 337
rect 702 335 716 337
rect 654 324 658 334
rect 664 333 668 335
rect 676 334 716 335
rect 664 331 665 333
rect 667 331 668 333
rect 664 330 668 331
rect 654 322 655 324
rect 657 322 658 324
rect 654 320 658 322
rect 661 326 668 330
rect 661 315 665 326
rect 704 321 708 326
rect 704 319 705 321
rect 707 319 708 321
rect 647 314 665 315
rect 647 312 649 314
rect 651 313 665 314
rect 651 312 676 313
rect 647 311 672 312
rect 661 310 672 311
rect 674 310 676 312
rect 661 309 676 310
rect 681 312 685 314
rect 681 310 682 312
rect 684 310 685 312
rect 681 305 685 310
rect 704 317 708 319
rect 712 323 716 334
rect 712 321 718 323
rect 712 319 715 321
rect 717 319 718 321
rect 712 317 718 319
rect 712 314 716 317
rect 696 310 716 314
rect 696 306 700 310
rect 660 304 682 305
rect 651 301 655 303
rect 660 302 662 304
rect 664 303 682 304
rect 684 303 685 305
rect 664 302 685 303
rect 690 305 700 306
rect 690 303 692 305
rect 694 303 700 305
rect 690 302 700 303
rect 751 338 755 342
rect 774 338 798 342
rect 738 337 778 338
rect 738 335 752 337
rect 754 335 778 337
rect 738 334 778 335
rect 738 323 742 334
rect 786 333 790 335
rect 794 334 800 338
rect 786 331 787 333
rect 789 331 790 333
rect 786 330 790 331
rect 786 326 793 330
rect 736 321 742 323
rect 736 319 737 321
rect 739 319 742 321
rect 736 317 742 319
rect 746 321 750 326
rect 746 319 747 321
rect 749 319 750 321
rect 746 317 750 319
rect 738 314 742 317
rect 738 310 758 314
rect 754 306 758 310
rect 789 315 793 326
rect 796 324 800 334
rect 796 322 797 324
rect 799 322 800 324
rect 796 320 800 322
rect 789 314 807 315
rect 769 312 773 314
rect 789 313 803 314
rect 769 310 770 312
rect 772 310 773 312
rect 754 305 764 306
rect 754 303 760 305
rect 762 303 764 305
rect 754 302 764 303
rect 769 305 773 310
rect 778 312 803 313
rect 805 312 807 314
rect 778 310 780 312
rect 782 311 807 312
rect 782 310 793 311
rect 778 309 793 310
rect 832 338 836 342
rect 832 334 847 338
rect 822 325 828 326
rect 843 321 847 334
rect 850 331 851 342
rect 843 319 844 321
rect 846 319 847 321
rect 843 313 847 319
rect 878 338 882 343
rect 887 343 893 352
rect 928 350 930 352
rect 932 350 934 352
rect 928 349 934 350
rect 963 350 965 352
rect 967 350 969 352
rect 887 341 889 343
rect 891 341 893 343
rect 963 345 969 350
rect 985 350 987 352
rect 989 350 991 352
rect 963 343 965 345
rect 967 343 969 345
rect 963 342 969 343
rect 976 344 980 346
rect 976 342 977 344
rect 979 342 980 344
rect 985 345 991 350
rect 985 343 987 345
rect 989 343 991 345
rect 985 342 991 343
rect 1017 350 1019 352
rect 1021 350 1023 352
rect 1017 345 1023 350
rect 1039 350 1041 352
rect 1043 350 1045 352
rect 1017 343 1019 345
rect 1021 343 1023 345
rect 1017 342 1023 343
rect 1028 344 1032 346
rect 1028 342 1029 344
rect 1031 342 1032 344
rect 1039 345 1045 350
rect 1074 350 1076 352
rect 1078 350 1080 352
rect 1074 349 1080 350
rect 1115 350 1117 352
rect 1119 350 1121 352
rect 1115 349 1121 350
rect 1039 343 1041 345
rect 1043 343 1045 345
rect 1039 342 1045 343
rect 1096 345 1113 346
rect 1096 343 1098 345
rect 1100 343 1113 345
rect 1096 342 1113 343
rect 887 340 893 341
rect 878 336 879 338
rect 881 337 882 338
rect 881 336 895 337
rect 878 333 895 336
rect 829 312 847 313
rect 829 310 831 312
rect 833 310 847 312
rect 829 309 847 310
rect 891 321 895 333
rect 891 319 892 321
rect 894 319 895 321
rect 891 314 895 319
rect 883 310 895 314
rect 883 306 887 310
rect 898 307 899 309
rect 769 303 770 305
rect 772 304 794 305
rect 772 303 790 304
rect 769 302 790 303
rect 792 302 794 304
rect 660 301 685 302
rect 769 301 794 302
rect 799 301 803 303
rect 867 305 887 306
rect 867 303 869 305
rect 871 303 887 305
rect 867 302 887 303
rect 933 338 957 342
rect 976 338 980 342
rect 931 334 937 338
rect 953 337 993 338
rect 953 335 977 337
rect 979 335 993 337
rect 931 324 935 334
rect 941 333 945 335
rect 953 334 993 335
rect 941 331 942 333
rect 944 331 945 333
rect 941 330 945 331
rect 931 322 932 324
rect 934 322 935 324
rect 931 320 935 322
rect 938 326 945 330
rect 938 315 942 326
rect 981 321 985 326
rect 981 319 982 321
rect 984 319 985 321
rect 924 314 942 315
rect 924 312 926 314
rect 928 313 942 314
rect 928 312 953 313
rect 924 311 949 312
rect 938 310 949 311
rect 951 310 953 312
rect 938 309 953 310
rect 958 312 962 314
rect 958 310 959 312
rect 961 310 962 312
rect 958 305 962 310
rect 981 317 985 319
rect 989 323 993 334
rect 989 321 995 323
rect 989 319 992 321
rect 994 319 995 321
rect 989 317 995 319
rect 989 314 993 317
rect 973 310 993 314
rect 973 306 977 310
rect 937 304 959 305
rect 928 301 932 303
rect 937 302 939 304
rect 941 303 959 304
rect 961 303 962 305
rect 941 302 962 303
rect 967 305 977 306
rect 967 303 969 305
rect 971 303 977 305
rect 967 302 977 303
rect 1028 338 1032 342
rect 1051 338 1075 342
rect 1015 337 1055 338
rect 1015 335 1029 337
rect 1031 335 1055 337
rect 1015 334 1055 335
rect 1015 323 1019 334
rect 1063 333 1067 335
rect 1071 334 1077 338
rect 1063 331 1064 333
rect 1066 331 1067 333
rect 1063 330 1067 331
rect 1063 326 1070 330
rect 1013 321 1019 323
rect 1013 319 1014 321
rect 1016 319 1019 321
rect 1013 317 1019 319
rect 1023 321 1027 326
rect 1023 319 1024 321
rect 1026 319 1027 321
rect 1023 317 1027 319
rect 1015 314 1019 317
rect 1015 310 1035 314
rect 1031 306 1035 310
rect 1066 315 1070 326
rect 1073 324 1077 334
rect 1073 322 1074 324
rect 1076 322 1077 324
rect 1073 320 1077 322
rect 1066 314 1084 315
rect 1046 312 1050 314
rect 1066 313 1080 314
rect 1046 310 1047 312
rect 1049 310 1050 312
rect 1031 305 1041 306
rect 1031 303 1037 305
rect 1039 303 1041 305
rect 1031 302 1041 303
rect 1046 305 1050 310
rect 1055 312 1080 313
rect 1082 312 1084 314
rect 1055 310 1057 312
rect 1059 311 1084 312
rect 1059 310 1070 311
rect 1055 309 1070 310
rect 1109 338 1113 342
rect 1109 334 1124 338
rect 1099 325 1105 326
rect 1120 321 1124 334
rect 1127 331 1128 342
rect 1120 319 1121 321
rect 1123 319 1124 321
rect 1120 313 1124 319
rect 1106 312 1124 313
rect 1106 310 1108 312
rect 1110 310 1124 312
rect 1106 309 1124 310
rect 1046 303 1047 305
rect 1049 304 1071 305
rect 1049 303 1067 304
rect 1046 302 1067 303
rect 1069 302 1071 304
rect 937 301 962 302
rect 1046 301 1071 302
rect 1076 301 1080 303
rect -204 299 -203 301
rect -201 299 -200 301
rect -56 299 -55 301
rect -53 299 -52 301
rect -204 296 -200 299
rect -148 298 -142 299
rect -148 296 -146 298
rect -144 296 -142 298
rect -114 298 -108 299
rect -114 296 -112 298
rect -110 296 -108 298
rect -56 296 -52 299
rect -36 299 -30 300
rect -36 297 -34 299
rect -32 297 -30 299
rect -36 296 -30 297
rect -17 299 -11 300
rect -17 297 -15 299
rect -13 297 -11 299
rect -17 296 -11 297
rect 98 299 99 301
rect 101 299 102 301
rect 246 299 247 301
rect 249 299 250 301
rect 98 296 102 299
rect 154 298 160 299
rect 154 296 156 298
rect 158 296 160 298
rect 188 298 194 299
rect 188 296 190 298
rect 192 296 194 298
rect 246 296 250 299
rect 266 299 272 300
rect 266 297 268 299
rect 270 297 272 299
rect 266 296 272 297
rect 285 299 291 300
rect 285 297 287 299
rect 289 297 291 299
rect 285 296 291 297
rect 375 299 376 301
rect 378 299 379 301
rect 523 299 524 301
rect 526 299 527 301
rect 375 296 379 299
rect 431 298 437 299
rect 431 296 433 298
rect 435 296 437 298
rect 465 298 471 299
rect 465 296 467 298
rect 469 296 471 298
rect 523 296 527 299
rect 543 299 549 300
rect 543 297 545 299
rect 547 297 549 299
rect 543 296 549 297
rect 562 299 568 300
rect 562 297 564 299
rect 566 297 568 299
rect 562 296 568 297
rect 651 299 652 301
rect 654 299 655 301
rect 799 299 800 301
rect 802 299 803 301
rect 651 296 655 299
rect 707 298 713 299
rect 707 296 709 298
rect 711 296 713 298
rect 741 298 747 299
rect 741 296 743 298
rect 745 296 747 298
rect 799 296 803 299
rect 819 299 825 300
rect 819 297 821 299
rect 823 297 825 299
rect 819 296 825 297
rect 838 299 844 300
rect 838 297 840 299
rect 842 297 844 299
rect 838 296 844 297
rect 928 299 929 301
rect 931 299 932 301
rect 1076 299 1077 301
rect 1079 299 1080 301
rect 928 296 932 299
rect 984 298 990 299
rect 984 296 986 298
rect 988 296 990 298
rect 1018 298 1024 299
rect 1018 296 1020 298
rect 1022 296 1024 298
rect 1076 296 1080 299
rect 1096 299 1102 300
rect 1096 297 1098 299
rect 1100 297 1102 299
rect 1096 296 1102 297
rect 1115 299 1121 300
rect 1115 297 1117 299
rect 1119 297 1121 299
rect 1115 296 1121 297
rect -269 274 -263 280
rect -204 277 -200 280
rect -148 278 -146 280
rect -144 278 -142 280
rect -148 277 -142 278
rect -114 278 -112 280
rect -110 278 -108 280
rect -114 277 -108 278
rect -56 277 -52 280
rect -204 275 -203 277
rect -201 275 -200 277
rect -56 275 -55 277
rect -53 275 -52 277
rect -36 279 -30 280
rect -36 277 -34 279
rect -32 277 -30 279
rect -36 276 -30 277
rect -17 279 -11 280
rect -17 277 -15 279
rect -13 277 -11 279
rect -17 276 -11 277
rect 98 277 102 280
rect 154 278 156 280
rect 158 278 160 280
rect 154 277 160 278
rect 188 278 190 280
rect 192 278 194 280
rect 188 277 194 278
rect 246 277 250 280
rect 98 275 99 277
rect 101 275 102 277
rect 246 275 247 277
rect 249 275 250 277
rect 266 279 272 280
rect 266 277 268 279
rect 270 277 272 279
rect 266 276 272 277
rect 285 279 291 280
rect 285 277 287 279
rect 289 277 291 279
rect 285 276 291 277
rect 375 277 379 280
rect 431 278 433 280
rect 435 278 437 280
rect 431 277 437 278
rect 465 278 467 280
rect 469 278 471 280
rect 465 277 471 278
rect 523 277 527 280
rect 375 275 376 277
rect 378 275 379 277
rect 523 275 524 277
rect 526 275 527 277
rect 543 279 549 280
rect 543 277 545 279
rect 547 277 549 279
rect 543 276 549 277
rect 562 279 568 280
rect 562 277 564 279
rect 566 277 568 279
rect 562 276 568 277
rect 651 277 655 280
rect 707 278 709 280
rect 711 278 713 280
rect 707 277 713 278
rect 741 278 743 280
rect 745 278 747 280
rect 741 277 747 278
rect 799 277 803 280
rect 651 275 652 277
rect 654 275 655 277
rect 799 275 800 277
rect 802 275 803 277
rect 819 279 825 280
rect 819 277 821 279
rect 823 277 825 279
rect 819 276 825 277
rect 838 279 844 280
rect 838 277 840 279
rect 842 277 844 279
rect 838 276 844 277
rect 928 277 932 280
rect 984 278 986 280
rect 988 278 990 280
rect 984 277 990 278
rect 1018 278 1020 280
rect 1022 278 1024 280
rect 1018 277 1024 278
rect 1076 277 1080 280
rect 928 275 929 277
rect 931 275 932 277
rect 1076 275 1077 277
rect 1079 275 1080 277
rect 1096 279 1102 280
rect 1096 277 1098 279
rect 1100 277 1102 279
rect 1096 276 1102 277
rect 1115 279 1121 280
rect 1115 277 1117 279
rect 1119 277 1121 279
rect 1115 276 1121 277
rect -269 272 -267 274
rect -265 272 -263 274
rect -269 271 -263 272
rect -256 271 -252 273
rect -256 269 -255 271
rect -253 269 -252 271
rect -282 266 -278 268
rect -282 264 -281 266
rect -279 264 -278 266
rect -282 258 -278 264
rect -256 266 -252 269
rect -256 262 -232 266
rect -282 254 -271 258
rect -275 248 -271 254
rect -236 258 -232 262
rect -256 257 -240 258
rect -256 255 -244 257
rect -242 255 -240 257
rect -256 254 -240 255
rect -236 256 -231 258
rect -236 254 -234 256
rect -232 254 -231 256
rect -256 248 -252 254
rect -236 252 -231 254
rect -236 250 -232 252
rect -275 247 -252 248
rect -275 245 -273 247
rect -271 245 -252 247
rect -275 244 -252 245
rect -264 233 -260 235
rect -264 231 -263 233
rect -261 231 -260 233
rect -264 226 -260 231
rect -256 233 -252 244
rect -248 247 -232 250
rect -248 245 -247 247
rect -245 246 -232 247
rect -245 245 -244 246
rect -248 240 -244 245
rect -248 238 -247 240
rect -245 238 -244 240
rect -248 236 -244 238
rect -204 273 -200 275
rect -195 274 -170 275
rect -86 274 -61 275
rect -195 272 -193 274
rect -191 273 -170 274
rect -191 272 -173 273
rect -195 271 -173 272
rect -171 271 -170 273
rect -194 266 -179 267
rect -194 265 -183 266
rect -208 264 -183 265
rect -181 264 -179 266
rect -208 262 -206 264
rect -204 263 -179 264
rect -174 266 -170 271
rect -165 273 -155 274
rect -165 271 -163 273
rect -161 271 -155 273
rect -165 270 -155 271
rect -174 264 -173 266
rect -171 264 -170 266
rect -204 262 -190 263
rect -174 262 -170 264
rect -208 261 -190 262
rect -201 254 -197 256
rect -201 252 -200 254
rect -198 252 -197 254
rect -201 242 -197 252
rect -194 250 -190 261
rect -159 266 -155 270
rect -159 262 -139 266
rect -143 259 -139 262
rect -151 257 -147 259
rect -151 255 -150 257
rect -148 255 -147 257
rect -151 250 -147 255
rect -143 257 -137 259
rect -143 255 -140 257
rect -138 255 -137 257
rect -143 253 -137 255
rect -194 246 -187 250
rect -191 245 -187 246
rect -191 243 -190 245
rect -188 243 -187 245
rect -201 238 -195 242
rect -191 241 -187 243
rect -143 242 -139 253
rect -179 241 -139 242
rect -179 239 -155 241
rect -153 239 -139 241
rect -179 238 -139 239
rect -199 234 -175 238
rect -156 234 -152 238
rect -101 273 -91 274
rect -101 271 -95 273
rect -93 271 -91 273
rect -101 270 -91 271
rect -86 273 -65 274
rect -86 271 -85 273
rect -83 272 -65 273
rect -63 272 -61 274
rect -56 273 -52 275
rect -83 271 -61 272
rect -101 266 -97 270
rect -117 262 -97 266
rect -117 259 -113 262
rect -119 257 -113 259
rect -119 255 -118 257
rect -116 255 -113 257
rect -119 253 -113 255
rect -117 242 -113 253
rect -109 257 -105 259
rect -86 266 -82 271
rect 7 273 27 274
rect 7 271 9 273
rect 11 271 27 273
rect 7 270 27 271
rect -86 264 -85 266
rect -83 264 -82 266
rect -86 262 -82 264
rect -77 266 -62 267
rect -77 264 -75 266
rect -73 265 -62 266
rect -73 264 -48 265
rect -77 263 -52 264
rect -66 262 -52 263
rect -50 262 -48 264
rect -66 261 -48 262
rect -109 255 -108 257
rect -106 255 -105 257
rect -109 250 -105 255
rect -66 250 -62 261
rect -69 246 -62 250
rect -59 254 -55 256
rect -59 252 -58 254
rect -56 252 -55 254
rect -69 245 -65 246
rect -69 243 -68 245
rect -66 243 -65 245
rect -117 241 -77 242
rect -69 241 -65 243
rect -59 242 -55 252
rect -26 266 -8 267
rect -26 264 -24 266
rect -22 264 -8 266
rect -26 263 -8 264
rect -12 257 -8 263
rect -12 255 -11 257
rect -9 255 -8 257
rect -33 250 -27 251
rect -117 239 -103 241
rect -101 239 -77 241
rect -117 238 -77 239
rect -61 238 -55 242
rect -104 234 -100 238
rect -81 234 -57 238
rect -12 242 -8 255
rect 23 266 27 270
rect 47 273 67 274
rect 47 271 49 273
rect 51 271 67 273
rect 47 270 67 271
rect 38 267 39 269
rect 23 262 35 266
rect 31 257 35 262
rect 31 255 32 257
rect 34 255 35 257
rect -23 238 -8 242
rect -23 234 -19 238
rect -5 234 -4 245
rect 31 243 35 255
rect 63 266 67 270
rect 78 267 79 269
rect 63 262 75 266
rect 71 257 75 262
rect 71 255 72 257
rect 74 255 75 257
rect 18 240 35 243
rect 18 238 19 240
rect 21 239 35 240
rect 21 238 22 239
rect -169 233 -163 234
rect -256 232 -223 233
rect -256 230 -227 232
rect -225 230 -223 232
rect -256 229 -223 230
rect -169 231 -167 233
rect -165 231 -163 233
rect -264 224 -263 226
rect -261 224 -260 226
rect -204 226 -198 227
rect -204 224 -202 226
rect -200 224 -198 226
rect -169 226 -163 231
rect -156 232 -155 234
rect -153 232 -152 234
rect -156 230 -152 232
rect -147 233 -141 234
rect -147 231 -145 233
rect -143 231 -141 233
rect -169 224 -167 226
rect -165 224 -163 226
rect -147 226 -141 231
rect -147 224 -145 226
rect -143 224 -141 226
rect -115 233 -109 234
rect -115 231 -113 233
rect -111 231 -109 233
rect -115 226 -109 231
rect -104 232 -103 234
rect -101 232 -100 234
rect -104 230 -100 232
rect -93 233 -87 234
rect -93 231 -91 233
rect -89 231 -87 233
rect -115 224 -113 226
rect -111 224 -109 226
rect -93 226 -87 231
rect -36 233 -19 234
rect -36 231 -34 233
rect -32 231 -19 233
rect -36 230 -19 231
rect 7 233 13 234
rect 7 231 9 233
rect 11 231 13 233
rect -93 224 -91 226
rect -89 224 -87 226
rect -58 226 -52 227
rect -58 224 -56 226
rect -54 224 -52 226
rect -17 226 -11 227
rect -17 224 -15 226
rect -13 224 -11 226
rect 7 224 13 231
rect 18 233 22 238
rect 71 243 75 255
rect 58 240 75 243
rect 58 238 59 240
rect 61 239 75 240
rect 61 238 62 239
rect 18 231 19 233
rect 21 231 22 233
rect 18 229 22 231
rect 27 235 33 236
rect 27 233 29 235
rect 31 233 33 235
rect 27 224 33 233
rect 47 233 53 234
rect 47 231 49 233
rect 51 231 53 233
rect 47 224 53 231
rect 58 233 62 238
rect 98 273 102 275
rect 107 274 132 275
rect 216 274 241 275
rect 107 272 109 274
rect 111 273 132 274
rect 111 272 129 273
rect 107 271 129 272
rect 131 271 132 273
rect 108 266 123 267
rect 108 265 119 266
rect 94 264 119 265
rect 121 264 123 266
rect 94 262 96 264
rect 98 263 123 264
rect 128 266 132 271
rect 137 273 147 274
rect 137 271 139 273
rect 141 271 147 273
rect 137 270 147 271
rect 128 264 129 266
rect 131 264 132 266
rect 98 262 112 263
rect 128 262 132 264
rect 94 261 112 262
rect 101 254 105 256
rect 101 252 102 254
rect 104 252 105 254
rect 101 242 105 252
rect 108 250 112 261
rect 143 266 147 270
rect 143 262 163 266
rect 159 259 163 262
rect 151 257 155 259
rect 151 255 152 257
rect 154 255 155 257
rect 151 250 155 255
rect 159 257 165 259
rect 159 255 162 257
rect 164 255 165 257
rect 159 253 165 255
rect 108 246 115 250
rect 111 245 115 246
rect 111 243 112 245
rect 114 243 115 245
rect 101 238 107 242
rect 111 241 115 243
rect 159 242 163 253
rect 123 241 163 242
rect 123 239 147 241
rect 149 239 163 241
rect 123 238 163 239
rect 58 231 59 233
rect 61 231 62 233
rect 58 229 62 231
rect 67 235 73 236
rect 67 233 69 235
rect 71 233 73 235
rect 103 234 127 238
rect 146 234 150 238
rect 201 273 211 274
rect 201 271 207 273
rect 209 271 211 273
rect 201 270 211 271
rect 216 273 237 274
rect 216 271 217 273
rect 219 272 237 273
rect 239 272 241 274
rect 246 273 250 275
rect 219 271 241 272
rect 201 266 205 270
rect 185 262 205 266
rect 185 259 189 262
rect 183 257 189 259
rect 183 255 184 257
rect 186 255 189 257
rect 183 253 189 255
rect 185 242 189 253
rect 193 257 197 259
rect 216 266 220 271
rect 314 273 334 274
rect 314 271 316 273
rect 318 271 334 273
rect 314 270 334 271
rect 216 264 217 266
rect 219 264 220 266
rect 216 262 220 264
rect 225 266 240 267
rect 225 264 227 266
rect 229 265 240 266
rect 229 264 254 265
rect 225 263 250 264
rect 236 262 250 263
rect 252 262 254 264
rect 236 261 254 262
rect 193 255 194 257
rect 196 255 197 257
rect 193 250 197 255
rect 236 250 240 261
rect 233 246 240 250
rect 243 254 247 256
rect 243 252 244 254
rect 246 252 247 254
rect 233 245 237 246
rect 233 243 234 245
rect 236 243 237 245
rect 185 241 225 242
rect 233 241 237 243
rect 243 242 247 252
rect 276 266 294 267
rect 276 264 278 266
rect 280 264 294 266
rect 276 263 294 264
rect 290 257 294 263
rect 290 255 291 257
rect 293 255 294 257
rect 269 250 275 251
rect 185 239 199 241
rect 201 239 225 241
rect 185 238 225 239
rect 241 238 247 242
rect 198 234 202 238
rect 221 234 245 238
rect 290 242 294 255
rect 279 238 294 242
rect 279 234 283 238
rect 297 234 298 245
rect 330 266 334 270
rect 345 267 346 269
rect 330 262 342 266
rect 338 257 342 262
rect 338 255 339 257
rect 341 255 342 257
rect 338 243 342 255
rect 325 240 342 243
rect 325 238 326 240
rect 328 239 342 240
rect 328 238 329 239
rect 67 224 73 233
rect 133 233 139 234
rect 133 231 135 233
rect 137 231 139 233
rect 98 226 104 227
rect 98 224 100 226
rect 102 224 104 226
rect 133 226 139 231
rect 146 232 147 234
rect 149 232 150 234
rect 146 230 150 232
rect 155 233 161 234
rect 155 231 157 233
rect 159 231 161 233
rect 133 224 135 226
rect 137 224 139 226
rect 155 226 161 231
rect 155 224 157 226
rect 159 224 161 226
rect 187 233 193 234
rect 187 231 189 233
rect 191 231 193 233
rect 187 226 193 231
rect 198 232 199 234
rect 201 232 202 234
rect 198 230 202 232
rect 209 233 215 234
rect 209 231 211 233
rect 213 231 215 233
rect 187 224 189 226
rect 191 224 193 226
rect 209 226 215 231
rect 266 233 283 234
rect 266 231 268 233
rect 270 231 283 233
rect 266 230 283 231
rect 314 233 320 234
rect 314 231 316 233
rect 318 231 320 233
rect 209 224 211 226
rect 213 224 215 226
rect 244 226 250 227
rect 244 224 246 226
rect 248 224 250 226
rect 285 226 291 227
rect 285 224 287 226
rect 289 224 291 226
rect 314 224 320 231
rect 325 233 329 238
rect 375 273 379 275
rect 384 274 409 275
rect 493 274 518 275
rect 384 272 386 274
rect 388 273 409 274
rect 388 272 406 273
rect 384 271 406 272
rect 408 271 409 273
rect 385 266 400 267
rect 385 265 396 266
rect 371 264 396 265
rect 398 264 400 266
rect 371 262 373 264
rect 375 263 400 264
rect 405 266 409 271
rect 414 273 424 274
rect 414 271 416 273
rect 418 271 424 273
rect 414 270 424 271
rect 405 264 406 266
rect 408 264 409 266
rect 375 262 389 263
rect 405 262 409 264
rect 371 261 389 262
rect 378 254 382 256
rect 378 252 379 254
rect 381 252 382 254
rect 378 242 382 252
rect 385 250 389 261
rect 420 266 424 270
rect 420 262 440 266
rect 436 259 440 262
rect 428 257 432 259
rect 428 255 429 257
rect 431 255 432 257
rect 428 250 432 255
rect 436 257 442 259
rect 436 255 439 257
rect 441 255 442 257
rect 436 253 442 255
rect 385 246 392 250
rect 388 245 392 246
rect 388 243 389 245
rect 391 243 392 245
rect 378 238 384 242
rect 388 241 392 243
rect 436 242 440 253
rect 400 241 440 242
rect 400 239 424 241
rect 426 239 440 241
rect 400 238 440 239
rect 325 231 326 233
rect 328 231 329 233
rect 325 229 329 231
rect 334 235 340 236
rect 334 233 336 235
rect 338 233 340 235
rect 380 234 404 238
rect 423 234 427 238
rect 478 273 488 274
rect 478 271 484 273
rect 486 271 488 273
rect 478 270 488 271
rect 493 273 514 274
rect 493 271 494 273
rect 496 272 514 273
rect 516 272 518 274
rect 523 273 527 275
rect 496 271 518 272
rect 478 266 482 270
rect 462 262 482 266
rect 462 259 466 262
rect 460 257 466 259
rect 460 255 461 257
rect 463 255 466 257
rect 460 253 466 255
rect 462 242 466 253
rect 470 257 474 259
rect 493 266 497 271
rect 591 273 611 274
rect 591 271 593 273
rect 595 271 611 273
rect 591 270 611 271
rect 493 264 494 266
rect 496 264 497 266
rect 493 262 497 264
rect 502 266 517 267
rect 502 264 504 266
rect 506 265 517 266
rect 506 264 531 265
rect 502 263 527 264
rect 513 262 527 263
rect 529 262 531 264
rect 513 261 531 262
rect 470 255 471 257
rect 473 255 474 257
rect 470 250 474 255
rect 513 250 517 261
rect 510 246 517 250
rect 520 254 524 256
rect 520 252 521 254
rect 523 252 524 254
rect 510 245 514 246
rect 510 243 511 245
rect 513 243 514 245
rect 462 241 502 242
rect 510 241 514 243
rect 520 242 524 252
rect 553 266 571 267
rect 553 264 555 266
rect 557 264 571 266
rect 553 263 571 264
rect 567 257 571 263
rect 567 255 568 257
rect 570 255 571 257
rect 546 250 552 251
rect 462 239 476 241
rect 478 239 502 241
rect 462 238 502 239
rect 518 238 524 242
rect 475 234 479 238
rect 498 234 522 238
rect 567 242 571 255
rect 556 238 571 242
rect 556 234 560 238
rect 574 234 575 245
rect 607 266 611 270
rect 622 267 623 269
rect 607 262 619 266
rect 615 257 619 262
rect 615 255 616 257
rect 618 255 619 257
rect 615 243 619 255
rect 602 240 619 243
rect 602 238 603 240
rect 605 239 619 240
rect 605 238 606 239
rect 334 224 340 233
rect 410 233 416 234
rect 410 231 412 233
rect 414 231 416 233
rect 375 226 381 227
rect 375 224 377 226
rect 379 224 381 226
rect 410 226 416 231
rect 423 232 424 234
rect 426 232 427 234
rect 423 230 427 232
rect 432 233 438 234
rect 432 231 434 233
rect 436 231 438 233
rect 410 224 412 226
rect 414 224 416 226
rect 432 226 438 231
rect 432 224 434 226
rect 436 224 438 226
rect 464 233 470 234
rect 464 231 466 233
rect 468 231 470 233
rect 464 226 470 231
rect 475 232 476 234
rect 478 232 479 234
rect 475 230 479 232
rect 486 233 492 234
rect 486 231 488 233
rect 490 231 492 233
rect 464 224 466 226
rect 468 224 470 226
rect 486 226 492 231
rect 543 233 560 234
rect 543 231 545 233
rect 547 231 560 233
rect 543 230 560 231
rect 591 233 597 234
rect 591 231 593 233
rect 595 231 597 233
rect 486 224 488 226
rect 490 224 492 226
rect 521 226 527 227
rect 521 224 523 226
rect 525 224 527 226
rect 562 226 568 227
rect 562 224 564 226
rect 566 224 568 226
rect 591 224 597 231
rect 602 233 606 238
rect 651 273 655 275
rect 660 274 685 275
rect 769 274 794 275
rect 660 272 662 274
rect 664 273 685 274
rect 664 272 682 273
rect 660 271 682 272
rect 684 271 685 273
rect 661 266 676 267
rect 661 265 672 266
rect 647 264 672 265
rect 674 264 676 266
rect 647 262 649 264
rect 651 263 676 264
rect 681 266 685 271
rect 690 273 700 274
rect 690 271 692 273
rect 694 271 700 273
rect 690 270 700 271
rect 681 264 682 266
rect 684 264 685 266
rect 651 262 665 263
rect 681 262 685 264
rect 647 261 665 262
rect 654 254 658 256
rect 654 252 655 254
rect 657 252 658 254
rect 654 242 658 252
rect 661 250 665 261
rect 696 266 700 270
rect 696 262 716 266
rect 712 259 716 262
rect 704 257 708 259
rect 704 255 705 257
rect 707 255 708 257
rect 704 250 708 255
rect 712 257 718 259
rect 712 255 715 257
rect 717 255 718 257
rect 712 253 718 255
rect 661 246 668 250
rect 664 245 668 246
rect 664 243 665 245
rect 667 243 668 245
rect 654 238 660 242
rect 664 241 668 243
rect 712 242 716 253
rect 676 241 716 242
rect 676 239 700 241
rect 702 239 716 241
rect 676 238 716 239
rect 602 231 603 233
rect 605 231 606 233
rect 602 229 606 231
rect 611 235 617 236
rect 611 233 613 235
rect 615 233 617 235
rect 656 234 680 238
rect 699 234 703 238
rect 754 273 764 274
rect 754 271 760 273
rect 762 271 764 273
rect 754 270 764 271
rect 769 273 790 274
rect 769 271 770 273
rect 772 272 790 273
rect 792 272 794 274
rect 799 273 803 275
rect 772 271 794 272
rect 754 266 758 270
rect 738 262 758 266
rect 738 259 742 262
rect 736 257 742 259
rect 736 255 737 257
rect 739 255 742 257
rect 736 253 742 255
rect 738 242 742 253
rect 746 257 750 259
rect 769 266 773 271
rect 867 273 887 274
rect 867 271 869 273
rect 871 271 887 273
rect 867 270 887 271
rect 769 264 770 266
rect 772 264 773 266
rect 769 262 773 264
rect 778 266 793 267
rect 778 264 780 266
rect 782 265 793 266
rect 782 264 807 265
rect 778 263 803 264
rect 789 262 803 263
rect 805 262 807 264
rect 789 261 807 262
rect 746 255 747 257
rect 749 255 750 257
rect 746 250 750 255
rect 789 250 793 261
rect 786 246 793 250
rect 796 254 800 256
rect 796 252 797 254
rect 799 252 800 254
rect 786 245 790 246
rect 786 243 787 245
rect 789 243 790 245
rect 738 241 778 242
rect 786 241 790 243
rect 796 242 800 252
rect 829 266 847 267
rect 829 264 831 266
rect 833 264 847 266
rect 829 263 847 264
rect 843 257 847 263
rect 843 255 844 257
rect 846 255 847 257
rect 822 250 828 251
rect 738 239 752 241
rect 754 239 778 241
rect 738 238 778 239
rect 794 238 800 242
rect 751 234 755 238
rect 774 234 798 238
rect 843 242 847 255
rect 832 238 847 242
rect 832 234 836 238
rect 850 234 851 245
rect 883 266 887 270
rect 898 267 899 269
rect 883 262 895 266
rect 891 257 895 262
rect 891 255 892 257
rect 894 255 895 257
rect 891 243 895 255
rect 878 240 895 243
rect 878 238 879 240
rect 881 239 895 240
rect 881 238 882 239
rect 611 224 617 233
rect 686 233 692 234
rect 686 231 688 233
rect 690 231 692 233
rect 651 226 657 227
rect 651 224 653 226
rect 655 224 657 226
rect 686 226 692 231
rect 699 232 700 234
rect 702 232 703 234
rect 699 230 703 232
rect 708 233 714 234
rect 708 231 710 233
rect 712 231 714 233
rect 686 224 688 226
rect 690 224 692 226
rect 708 226 714 231
rect 708 224 710 226
rect 712 224 714 226
rect 740 233 746 234
rect 740 231 742 233
rect 744 231 746 233
rect 740 226 746 231
rect 751 232 752 234
rect 754 232 755 234
rect 751 230 755 232
rect 762 233 768 234
rect 762 231 764 233
rect 766 231 768 233
rect 740 224 742 226
rect 744 224 746 226
rect 762 226 768 231
rect 819 233 836 234
rect 819 231 821 233
rect 823 231 836 233
rect 819 230 836 231
rect 867 233 873 234
rect 867 231 869 233
rect 871 231 873 233
rect 762 224 764 226
rect 766 224 768 226
rect 797 226 803 227
rect 797 224 799 226
rect 801 224 803 226
rect 838 226 844 227
rect 838 224 840 226
rect 842 224 844 226
rect 867 224 873 231
rect 878 233 882 238
rect 928 273 932 275
rect 937 274 962 275
rect 1046 274 1071 275
rect 937 272 939 274
rect 941 273 962 274
rect 941 272 959 273
rect 937 271 959 272
rect 961 271 962 273
rect 938 266 953 267
rect 938 265 949 266
rect 924 264 949 265
rect 951 264 953 266
rect 924 262 926 264
rect 928 263 953 264
rect 958 266 962 271
rect 967 273 977 274
rect 967 271 969 273
rect 971 271 977 273
rect 967 270 977 271
rect 958 264 959 266
rect 961 264 962 266
rect 928 262 942 263
rect 958 262 962 264
rect 924 261 942 262
rect 931 254 935 256
rect 931 252 932 254
rect 934 252 935 254
rect 931 242 935 252
rect 938 250 942 261
rect 973 266 977 270
rect 973 262 993 266
rect 989 259 993 262
rect 981 257 985 259
rect 981 255 982 257
rect 984 255 985 257
rect 981 250 985 255
rect 989 257 995 259
rect 989 255 992 257
rect 994 255 995 257
rect 989 253 995 255
rect 938 246 945 250
rect 941 245 945 246
rect 941 243 942 245
rect 944 243 945 245
rect 931 238 937 242
rect 941 241 945 243
rect 989 242 993 253
rect 953 241 993 242
rect 953 239 977 241
rect 979 239 993 241
rect 953 238 993 239
rect 878 231 879 233
rect 881 231 882 233
rect 878 229 882 231
rect 887 235 893 236
rect 887 233 889 235
rect 891 233 893 235
rect 933 234 957 238
rect 976 234 980 238
rect 1031 273 1041 274
rect 1031 271 1037 273
rect 1039 271 1041 273
rect 1031 270 1041 271
rect 1046 273 1067 274
rect 1046 271 1047 273
rect 1049 272 1067 273
rect 1069 272 1071 274
rect 1076 273 1080 275
rect 1049 271 1071 272
rect 1031 266 1035 270
rect 1015 262 1035 266
rect 1015 259 1019 262
rect 1013 257 1019 259
rect 1013 255 1014 257
rect 1016 255 1019 257
rect 1013 253 1019 255
rect 1015 242 1019 253
rect 1023 257 1027 259
rect 1046 266 1050 271
rect 1046 264 1047 266
rect 1049 264 1050 266
rect 1046 262 1050 264
rect 1055 266 1070 267
rect 1055 264 1057 266
rect 1059 265 1070 266
rect 1059 264 1084 265
rect 1055 263 1080 264
rect 1066 262 1080 263
rect 1082 262 1084 264
rect 1066 261 1084 262
rect 1023 255 1024 257
rect 1026 255 1027 257
rect 1023 250 1027 255
rect 1066 250 1070 261
rect 1063 246 1070 250
rect 1073 254 1077 256
rect 1073 252 1074 254
rect 1076 252 1077 254
rect 1063 245 1067 246
rect 1063 243 1064 245
rect 1066 243 1067 245
rect 1015 241 1055 242
rect 1063 241 1067 243
rect 1073 242 1077 252
rect 1106 266 1124 267
rect 1106 264 1108 266
rect 1110 264 1124 266
rect 1106 263 1124 264
rect 1120 257 1124 263
rect 1120 255 1121 257
rect 1123 255 1124 257
rect 1099 250 1105 251
rect 1015 239 1029 241
rect 1031 239 1055 241
rect 1015 238 1055 239
rect 1071 238 1077 242
rect 1028 234 1032 238
rect 1051 234 1075 238
rect 1120 242 1124 255
rect 1109 238 1124 242
rect 1109 234 1113 238
rect 1127 234 1128 245
rect 887 224 893 233
rect 963 233 969 234
rect 963 231 965 233
rect 967 231 969 233
rect 928 226 934 227
rect 928 224 930 226
rect 932 224 934 226
rect 963 226 969 231
rect 976 232 977 234
rect 979 232 980 234
rect 976 230 980 232
rect 985 233 991 234
rect 985 231 987 233
rect 989 231 991 233
rect 963 224 965 226
rect 967 224 969 226
rect 985 226 991 231
rect 985 224 987 226
rect 989 224 991 226
rect 1017 233 1023 234
rect 1017 231 1019 233
rect 1021 231 1023 233
rect 1017 226 1023 231
rect 1028 232 1029 234
rect 1031 232 1032 234
rect 1028 230 1032 232
rect 1039 233 1045 234
rect 1039 231 1041 233
rect 1043 231 1045 233
rect 1017 224 1019 226
rect 1021 224 1023 226
rect 1039 226 1045 231
rect 1096 233 1113 234
rect 1096 231 1098 233
rect 1100 231 1113 233
rect 1096 230 1113 231
rect 1039 224 1041 226
rect 1043 224 1045 226
rect 1074 226 1080 227
rect 1074 224 1076 226
rect 1078 224 1080 226
rect 1115 226 1121 227
rect 1115 224 1117 226
rect 1119 224 1121 226
rect -264 206 -263 208
rect -261 206 -260 208
rect -264 201 -260 206
rect -204 206 -202 208
rect -200 206 -198 208
rect -204 205 -198 206
rect -169 206 -167 208
rect -165 206 -163 208
rect -264 199 -263 201
rect -261 199 -260 201
rect -264 197 -260 199
rect -256 202 -223 203
rect -256 200 -227 202
rect -225 200 -223 202
rect -256 199 -223 200
rect -169 201 -163 206
rect -147 206 -145 208
rect -143 206 -141 208
rect -169 199 -167 201
rect -165 199 -163 201
rect -256 188 -252 199
rect -169 198 -163 199
rect -156 200 -152 202
rect -156 198 -155 200
rect -153 198 -152 200
rect -147 201 -141 206
rect -147 199 -145 201
rect -143 199 -141 201
rect -147 198 -141 199
rect -115 206 -113 208
rect -111 206 -109 208
rect -115 201 -109 206
rect -93 206 -91 208
rect -89 206 -87 208
rect -115 199 -113 201
rect -111 199 -109 201
rect -115 198 -109 199
rect -104 200 -100 202
rect -104 198 -103 200
rect -101 198 -100 200
rect -93 201 -87 206
rect -58 206 -56 208
rect -54 206 -52 208
rect -58 205 -52 206
rect -17 206 -15 208
rect -13 206 -11 208
rect -17 205 -11 206
rect -93 199 -91 201
rect -89 199 -87 201
rect -93 198 -87 199
rect -36 201 -19 202
rect -36 199 -34 201
rect -32 199 -19 201
rect -36 198 -19 199
rect 7 201 13 208
rect 7 199 9 201
rect 11 199 13 201
rect 7 198 13 199
rect 18 201 22 203
rect 18 199 19 201
rect 21 199 22 201
rect -275 187 -252 188
rect -275 185 -273 187
rect -271 185 -252 187
rect -275 184 -252 185
rect -275 178 -271 184
rect -282 174 -271 178
rect -282 168 -278 174
rect -256 178 -252 184
rect -248 194 -244 196
rect -248 192 -247 194
rect -245 192 -244 194
rect -248 187 -244 192
rect -248 185 -247 187
rect -245 186 -244 187
rect -245 185 -232 186
rect -248 182 -232 185
rect -236 180 -232 182
rect -236 178 -231 180
rect -256 177 -240 178
rect -256 175 -244 177
rect -242 175 -240 177
rect -256 174 -240 175
rect -236 176 -234 178
rect -232 176 -231 178
rect -236 174 -231 176
rect -282 166 -281 168
rect -279 166 -278 168
rect -282 164 -278 166
rect -236 170 -232 174
rect -256 166 -232 170
rect -256 163 -252 166
rect -256 161 -255 163
rect -253 161 -252 163
rect -269 160 -263 161
rect -269 158 -267 160
rect -265 158 -263 160
rect -256 159 -252 161
rect -199 194 -175 198
rect -156 194 -152 198
rect -201 190 -195 194
rect -179 193 -139 194
rect -179 191 -155 193
rect -153 191 -139 193
rect -201 180 -197 190
rect -191 189 -187 191
rect -179 190 -139 191
rect -191 187 -190 189
rect -188 187 -187 189
rect -191 186 -187 187
rect -201 178 -200 180
rect -198 178 -197 180
rect -201 176 -197 178
rect -194 182 -187 186
rect -194 171 -190 182
rect -151 177 -147 182
rect -151 175 -150 177
rect -148 175 -147 177
rect -208 170 -190 171
rect -208 168 -206 170
rect -204 169 -190 170
rect -204 168 -179 169
rect -208 167 -183 168
rect -194 166 -183 167
rect -181 166 -179 168
rect -194 165 -179 166
rect -174 168 -170 170
rect -174 166 -173 168
rect -171 166 -170 168
rect -174 161 -170 166
rect -151 173 -147 175
rect -143 179 -139 190
rect -143 177 -137 179
rect -143 175 -140 177
rect -138 175 -137 177
rect -143 173 -137 175
rect -143 170 -139 173
rect -159 166 -139 170
rect -159 162 -155 166
rect -195 160 -173 161
rect -269 152 -263 158
rect -204 157 -200 159
rect -195 158 -193 160
rect -191 159 -173 160
rect -171 159 -170 161
rect -191 158 -170 159
rect -165 161 -155 162
rect -165 159 -163 161
rect -161 159 -155 161
rect -165 158 -155 159
rect -104 194 -100 198
rect -81 194 -57 198
rect -117 193 -77 194
rect -117 191 -103 193
rect -101 191 -77 193
rect -117 190 -77 191
rect -117 179 -113 190
rect -69 189 -65 191
rect -61 190 -55 194
rect -69 187 -68 189
rect -66 187 -65 189
rect -69 186 -65 187
rect -69 182 -62 186
rect -119 177 -113 179
rect -119 175 -118 177
rect -116 175 -113 177
rect -119 173 -113 175
rect -109 177 -105 182
rect -109 175 -108 177
rect -106 175 -105 177
rect -109 173 -105 175
rect -117 170 -113 173
rect -117 166 -97 170
rect -101 162 -97 166
rect -66 171 -62 182
rect -59 180 -55 190
rect -59 178 -58 180
rect -56 178 -55 180
rect -59 176 -55 178
rect -66 170 -48 171
rect -86 168 -82 170
rect -66 169 -52 170
rect -86 166 -85 168
rect -83 166 -82 168
rect -101 161 -91 162
rect -101 159 -95 161
rect -93 159 -91 161
rect -101 158 -91 159
rect -86 161 -82 166
rect -77 168 -52 169
rect -50 168 -48 170
rect -77 166 -75 168
rect -73 167 -48 168
rect -23 194 -19 198
rect -23 190 -8 194
rect -33 181 -27 182
rect -73 166 -62 167
rect -77 165 -62 166
rect -12 177 -8 190
rect -5 187 -4 198
rect -12 175 -11 177
rect -9 175 -8 177
rect -12 169 -8 175
rect 18 194 22 199
rect 27 199 33 208
rect 47 201 53 208
rect 47 199 49 201
rect 51 199 53 201
rect 27 197 29 199
rect 31 197 33 199
rect 27 196 33 197
rect 47 198 53 199
rect 58 201 62 203
rect 58 199 59 201
rect 61 199 62 201
rect 18 192 19 194
rect 21 193 22 194
rect 21 192 35 193
rect 18 189 35 192
rect -26 168 -8 169
rect -26 166 -24 168
rect -22 166 -8 168
rect -26 165 -8 166
rect 31 177 35 189
rect 58 194 62 199
rect 67 199 73 208
rect 98 206 100 208
rect 102 206 104 208
rect 98 205 104 206
rect 133 206 135 208
rect 137 206 139 208
rect 67 197 69 199
rect 71 197 73 199
rect 133 201 139 206
rect 155 206 157 208
rect 159 206 161 208
rect 133 199 135 201
rect 137 199 139 201
rect 133 198 139 199
rect 146 200 150 202
rect 146 198 147 200
rect 149 198 150 200
rect 155 201 161 206
rect 155 199 157 201
rect 159 199 161 201
rect 155 198 161 199
rect 187 206 189 208
rect 191 206 193 208
rect 187 201 193 206
rect 209 206 211 208
rect 213 206 215 208
rect 187 199 189 201
rect 191 199 193 201
rect 187 198 193 199
rect 198 200 202 202
rect 198 198 199 200
rect 201 198 202 200
rect 209 201 215 206
rect 244 206 246 208
rect 248 206 250 208
rect 244 205 250 206
rect 285 206 287 208
rect 289 206 291 208
rect 285 205 291 206
rect 209 199 211 201
rect 213 199 215 201
rect 209 198 215 199
rect 266 201 283 202
rect 266 199 268 201
rect 270 199 283 201
rect 266 198 283 199
rect 314 201 320 208
rect 314 199 316 201
rect 318 199 320 201
rect 314 198 320 199
rect 325 201 329 203
rect 325 199 326 201
rect 328 199 329 201
rect 67 196 73 197
rect 58 192 59 194
rect 61 193 62 194
rect 61 192 75 193
rect 58 189 75 192
rect 31 175 32 177
rect 34 175 35 177
rect 31 170 35 175
rect 23 166 35 170
rect 23 162 27 166
rect 38 163 39 165
rect 71 177 75 189
rect 71 175 72 177
rect 74 175 75 177
rect 71 170 75 175
rect 63 166 75 170
rect -86 159 -85 161
rect -83 160 -61 161
rect -83 159 -65 160
rect -86 158 -65 159
rect -63 158 -61 160
rect -195 157 -170 158
rect -86 157 -61 158
rect -56 157 -52 159
rect 7 161 27 162
rect 7 159 9 161
rect 11 159 27 161
rect 7 158 27 159
rect 63 162 67 166
rect 78 163 79 165
rect 47 161 67 162
rect 47 159 49 161
rect 51 159 67 161
rect 47 158 67 159
rect 103 194 127 198
rect 146 194 150 198
rect 101 190 107 194
rect 123 193 163 194
rect 123 191 147 193
rect 149 191 163 193
rect 101 180 105 190
rect 111 189 115 191
rect 123 190 163 191
rect 111 187 112 189
rect 114 187 115 189
rect 111 186 115 187
rect 101 178 102 180
rect 104 178 105 180
rect 101 176 105 178
rect 108 182 115 186
rect 108 171 112 182
rect 151 177 155 182
rect 151 175 152 177
rect 154 175 155 177
rect 94 170 112 171
rect 94 168 96 170
rect 98 169 112 170
rect 98 168 123 169
rect 94 167 119 168
rect 108 166 119 167
rect 121 166 123 168
rect 108 165 123 166
rect 128 168 132 170
rect 128 166 129 168
rect 131 166 132 168
rect 128 161 132 166
rect 151 173 155 175
rect 159 179 163 190
rect 159 177 165 179
rect 159 175 162 177
rect 164 175 165 177
rect 159 173 165 175
rect 159 170 163 173
rect 143 166 163 170
rect 143 162 147 166
rect 107 160 129 161
rect 98 157 102 159
rect 107 158 109 160
rect 111 159 129 160
rect 131 159 132 161
rect 111 158 132 159
rect 137 161 147 162
rect 137 159 139 161
rect 141 159 147 161
rect 137 158 147 159
rect 198 194 202 198
rect 221 194 245 198
rect 185 193 225 194
rect 185 191 199 193
rect 201 191 225 193
rect 185 190 225 191
rect 185 179 189 190
rect 233 189 237 191
rect 241 190 247 194
rect 233 187 234 189
rect 236 187 237 189
rect 233 186 237 187
rect 233 182 240 186
rect 183 177 189 179
rect 183 175 184 177
rect 186 175 189 177
rect 183 173 189 175
rect 193 177 197 182
rect 193 175 194 177
rect 196 175 197 177
rect 193 173 197 175
rect 185 170 189 173
rect 185 166 205 170
rect 201 162 205 166
rect 236 171 240 182
rect 243 180 247 190
rect 243 178 244 180
rect 246 178 247 180
rect 243 176 247 178
rect 236 170 254 171
rect 216 168 220 170
rect 236 169 250 170
rect 216 166 217 168
rect 219 166 220 168
rect 201 161 211 162
rect 201 159 207 161
rect 209 159 211 161
rect 201 158 211 159
rect 216 161 220 166
rect 225 168 250 169
rect 252 168 254 170
rect 225 166 227 168
rect 229 167 254 168
rect 229 166 240 167
rect 225 165 240 166
rect 279 194 283 198
rect 279 190 294 194
rect 269 181 275 182
rect 290 177 294 190
rect 297 187 298 198
rect 290 175 291 177
rect 293 175 294 177
rect 290 169 294 175
rect 325 194 329 199
rect 334 199 340 208
rect 375 206 377 208
rect 379 206 381 208
rect 375 205 381 206
rect 410 206 412 208
rect 414 206 416 208
rect 334 197 336 199
rect 338 197 340 199
rect 410 201 416 206
rect 432 206 434 208
rect 436 206 438 208
rect 410 199 412 201
rect 414 199 416 201
rect 410 198 416 199
rect 423 200 427 202
rect 423 198 424 200
rect 426 198 427 200
rect 432 201 438 206
rect 432 199 434 201
rect 436 199 438 201
rect 432 198 438 199
rect 464 206 466 208
rect 468 206 470 208
rect 464 201 470 206
rect 486 206 488 208
rect 490 206 492 208
rect 464 199 466 201
rect 468 199 470 201
rect 464 198 470 199
rect 475 200 479 202
rect 475 198 476 200
rect 478 198 479 200
rect 486 201 492 206
rect 521 206 523 208
rect 525 206 527 208
rect 521 205 527 206
rect 562 206 564 208
rect 566 206 568 208
rect 562 205 568 206
rect 486 199 488 201
rect 490 199 492 201
rect 486 198 492 199
rect 543 201 560 202
rect 543 199 545 201
rect 547 199 560 201
rect 543 198 560 199
rect 591 201 597 208
rect 591 199 593 201
rect 595 199 597 201
rect 591 198 597 199
rect 602 201 606 203
rect 602 199 603 201
rect 605 199 606 201
rect 334 196 340 197
rect 325 192 326 194
rect 328 193 329 194
rect 328 192 342 193
rect 325 189 342 192
rect 276 168 294 169
rect 276 166 278 168
rect 280 166 294 168
rect 276 165 294 166
rect 338 177 342 189
rect 338 175 339 177
rect 341 175 342 177
rect 338 170 342 175
rect 330 166 342 170
rect 330 162 334 166
rect 345 163 346 165
rect 216 159 217 161
rect 219 160 241 161
rect 219 159 237 160
rect 216 158 237 159
rect 239 158 241 160
rect 107 157 132 158
rect 216 157 241 158
rect 246 157 250 159
rect 314 161 334 162
rect 314 159 316 161
rect 318 159 334 161
rect 314 158 334 159
rect 380 194 404 198
rect 423 194 427 198
rect 378 190 384 194
rect 400 193 440 194
rect 400 191 424 193
rect 426 191 440 193
rect 378 180 382 190
rect 388 189 392 191
rect 400 190 440 191
rect 388 187 389 189
rect 391 187 392 189
rect 388 186 392 187
rect 378 178 379 180
rect 381 178 382 180
rect 378 176 382 178
rect 385 182 392 186
rect 385 171 389 182
rect 428 177 432 182
rect 428 175 429 177
rect 431 175 432 177
rect 371 170 389 171
rect 371 168 373 170
rect 375 169 389 170
rect 375 168 400 169
rect 371 167 396 168
rect 385 166 396 167
rect 398 166 400 168
rect 385 165 400 166
rect 405 168 409 170
rect 405 166 406 168
rect 408 166 409 168
rect 405 161 409 166
rect 428 173 432 175
rect 436 179 440 190
rect 436 177 442 179
rect 436 175 439 177
rect 441 175 442 177
rect 436 173 442 175
rect 436 170 440 173
rect 420 166 440 170
rect 420 162 424 166
rect 384 160 406 161
rect 375 157 379 159
rect 384 158 386 160
rect 388 159 406 160
rect 408 159 409 161
rect 388 158 409 159
rect 414 161 424 162
rect 414 159 416 161
rect 418 159 424 161
rect 414 158 424 159
rect 475 194 479 198
rect 498 194 522 198
rect 462 193 502 194
rect 462 191 476 193
rect 478 191 502 193
rect 462 190 502 191
rect 462 179 466 190
rect 510 189 514 191
rect 518 190 524 194
rect 510 187 511 189
rect 513 187 514 189
rect 510 186 514 187
rect 510 182 517 186
rect 460 177 466 179
rect 460 175 461 177
rect 463 175 466 177
rect 460 173 466 175
rect 470 177 474 182
rect 470 175 471 177
rect 473 175 474 177
rect 470 173 474 175
rect 462 170 466 173
rect 462 166 482 170
rect 478 162 482 166
rect 513 171 517 182
rect 520 180 524 190
rect 520 178 521 180
rect 523 178 524 180
rect 520 176 524 178
rect 513 170 531 171
rect 493 168 497 170
rect 513 169 527 170
rect 493 166 494 168
rect 496 166 497 168
rect 478 161 488 162
rect 478 159 484 161
rect 486 159 488 161
rect 478 158 488 159
rect 493 161 497 166
rect 502 168 527 169
rect 529 168 531 170
rect 502 166 504 168
rect 506 167 531 168
rect 506 166 517 167
rect 502 165 517 166
rect 556 194 560 198
rect 556 190 571 194
rect 546 181 552 182
rect 567 177 571 190
rect 574 187 575 198
rect 567 175 568 177
rect 570 175 571 177
rect 567 169 571 175
rect 602 194 606 199
rect 611 199 617 208
rect 651 206 653 208
rect 655 206 657 208
rect 651 205 657 206
rect 686 206 688 208
rect 690 206 692 208
rect 611 197 613 199
rect 615 197 617 199
rect 686 201 692 206
rect 708 206 710 208
rect 712 206 714 208
rect 686 199 688 201
rect 690 199 692 201
rect 686 198 692 199
rect 699 200 703 202
rect 699 198 700 200
rect 702 198 703 200
rect 708 201 714 206
rect 708 199 710 201
rect 712 199 714 201
rect 708 198 714 199
rect 740 206 742 208
rect 744 206 746 208
rect 740 201 746 206
rect 762 206 764 208
rect 766 206 768 208
rect 740 199 742 201
rect 744 199 746 201
rect 740 198 746 199
rect 751 200 755 202
rect 751 198 752 200
rect 754 198 755 200
rect 762 201 768 206
rect 797 206 799 208
rect 801 206 803 208
rect 797 205 803 206
rect 838 206 840 208
rect 842 206 844 208
rect 838 205 844 206
rect 762 199 764 201
rect 766 199 768 201
rect 762 198 768 199
rect 819 201 836 202
rect 819 199 821 201
rect 823 199 836 201
rect 819 198 836 199
rect 867 201 873 208
rect 867 199 869 201
rect 871 199 873 201
rect 867 198 873 199
rect 878 201 882 203
rect 878 199 879 201
rect 881 199 882 201
rect 611 196 617 197
rect 602 192 603 194
rect 605 193 606 194
rect 605 192 619 193
rect 602 189 619 192
rect 553 168 571 169
rect 553 166 555 168
rect 557 166 571 168
rect 553 165 571 166
rect 615 177 619 189
rect 615 175 616 177
rect 618 175 619 177
rect 615 170 619 175
rect 607 166 619 170
rect 607 162 611 166
rect 622 163 623 165
rect 493 159 494 161
rect 496 160 518 161
rect 496 159 514 160
rect 493 158 514 159
rect 516 158 518 160
rect 384 157 409 158
rect 493 157 518 158
rect 523 157 527 159
rect 591 161 611 162
rect 591 159 593 161
rect 595 159 611 161
rect 591 158 611 159
rect 656 194 680 198
rect 699 194 703 198
rect 654 190 660 194
rect 676 193 716 194
rect 676 191 700 193
rect 702 191 716 193
rect 654 180 658 190
rect 664 189 668 191
rect 676 190 716 191
rect 664 187 665 189
rect 667 187 668 189
rect 664 186 668 187
rect 654 178 655 180
rect 657 178 658 180
rect 654 176 658 178
rect 661 182 668 186
rect 661 171 665 182
rect 704 177 708 182
rect 704 175 705 177
rect 707 175 708 177
rect 647 170 665 171
rect 647 168 649 170
rect 651 169 665 170
rect 651 168 676 169
rect 647 167 672 168
rect 661 166 672 167
rect 674 166 676 168
rect 661 165 676 166
rect 681 168 685 170
rect 681 166 682 168
rect 684 166 685 168
rect 681 161 685 166
rect 704 173 708 175
rect 712 179 716 190
rect 712 177 718 179
rect 712 175 715 177
rect 717 175 718 177
rect 712 173 718 175
rect 712 170 716 173
rect 696 166 716 170
rect 696 162 700 166
rect 660 160 682 161
rect 651 157 655 159
rect 660 158 662 160
rect 664 159 682 160
rect 684 159 685 161
rect 664 158 685 159
rect 690 161 700 162
rect 690 159 692 161
rect 694 159 700 161
rect 690 158 700 159
rect 751 194 755 198
rect 774 194 798 198
rect 738 193 778 194
rect 738 191 752 193
rect 754 191 778 193
rect 738 190 778 191
rect 738 179 742 190
rect 786 189 790 191
rect 794 190 800 194
rect 786 187 787 189
rect 789 187 790 189
rect 786 186 790 187
rect 786 182 793 186
rect 736 177 742 179
rect 736 175 737 177
rect 739 175 742 177
rect 736 173 742 175
rect 746 177 750 182
rect 746 175 747 177
rect 749 175 750 177
rect 746 173 750 175
rect 738 170 742 173
rect 738 166 758 170
rect 754 162 758 166
rect 789 171 793 182
rect 796 180 800 190
rect 796 178 797 180
rect 799 178 800 180
rect 796 176 800 178
rect 789 170 807 171
rect 769 168 773 170
rect 789 169 803 170
rect 769 166 770 168
rect 772 166 773 168
rect 754 161 764 162
rect 754 159 760 161
rect 762 159 764 161
rect 754 158 764 159
rect 769 161 773 166
rect 778 168 803 169
rect 805 168 807 170
rect 778 166 780 168
rect 782 167 807 168
rect 782 166 793 167
rect 778 165 793 166
rect 832 194 836 198
rect 832 190 847 194
rect 822 181 828 182
rect 843 177 847 190
rect 850 187 851 198
rect 843 175 844 177
rect 846 175 847 177
rect 843 169 847 175
rect 878 194 882 199
rect 887 199 893 208
rect 928 206 930 208
rect 932 206 934 208
rect 928 205 934 206
rect 963 206 965 208
rect 967 206 969 208
rect 887 197 889 199
rect 891 197 893 199
rect 963 201 969 206
rect 985 206 987 208
rect 989 206 991 208
rect 963 199 965 201
rect 967 199 969 201
rect 963 198 969 199
rect 976 200 980 202
rect 976 198 977 200
rect 979 198 980 200
rect 985 201 991 206
rect 985 199 987 201
rect 989 199 991 201
rect 985 198 991 199
rect 1017 206 1019 208
rect 1021 206 1023 208
rect 1017 201 1023 206
rect 1039 206 1041 208
rect 1043 206 1045 208
rect 1017 199 1019 201
rect 1021 199 1023 201
rect 1017 198 1023 199
rect 1028 200 1032 202
rect 1028 198 1029 200
rect 1031 198 1032 200
rect 1039 201 1045 206
rect 1074 206 1076 208
rect 1078 206 1080 208
rect 1074 205 1080 206
rect 1115 206 1117 208
rect 1119 206 1121 208
rect 1115 205 1121 206
rect 1039 199 1041 201
rect 1043 199 1045 201
rect 1039 198 1045 199
rect 1096 201 1113 202
rect 1096 199 1098 201
rect 1100 199 1113 201
rect 1096 198 1113 199
rect 887 196 893 197
rect 878 192 879 194
rect 881 193 882 194
rect 881 192 895 193
rect 878 189 895 192
rect 829 168 847 169
rect 829 166 831 168
rect 833 166 847 168
rect 829 165 847 166
rect 891 177 895 189
rect 891 175 892 177
rect 894 175 895 177
rect 891 170 895 175
rect 883 166 895 170
rect 883 162 887 166
rect 898 163 899 165
rect 769 159 770 161
rect 772 160 794 161
rect 772 159 790 160
rect 769 158 790 159
rect 792 158 794 160
rect 660 157 685 158
rect 769 157 794 158
rect 799 157 803 159
rect 867 161 887 162
rect 867 159 869 161
rect 871 159 887 161
rect 867 158 887 159
rect 933 194 957 198
rect 976 194 980 198
rect 931 190 937 194
rect 953 193 993 194
rect 953 191 977 193
rect 979 191 993 193
rect 931 180 935 190
rect 941 189 945 191
rect 953 190 993 191
rect 941 187 942 189
rect 944 187 945 189
rect 941 186 945 187
rect 931 178 932 180
rect 934 178 935 180
rect 931 176 935 178
rect 938 182 945 186
rect 938 171 942 182
rect 981 177 985 182
rect 981 175 982 177
rect 984 175 985 177
rect 924 170 942 171
rect 924 168 926 170
rect 928 169 942 170
rect 928 168 953 169
rect 924 167 949 168
rect 938 166 949 167
rect 951 166 953 168
rect 938 165 953 166
rect 958 168 962 170
rect 958 166 959 168
rect 961 166 962 168
rect 958 161 962 166
rect 981 173 985 175
rect 989 179 993 190
rect 989 177 995 179
rect 989 175 992 177
rect 994 175 995 177
rect 989 173 995 175
rect 989 170 993 173
rect 973 166 993 170
rect 973 162 977 166
rect 937 160 959 161
rect 928 157 932 159
rect 937 158 939 160
rect 941 159 959 160
rect 961 159 962 161
rect 941 158 962 159
rect 967 161 977 162
rect 967 159 969 161
rect 971 159 977 161
rect 967 158 977 159
rect 1028 194 1032 198
rect 1051 194 1075 198
rect 1015 193 1055 194
rect 1015 191 1029 193
rect 1031 191 1055 193
rect 1015 190 1055 191
rect 1015 179 1019 190
rect 1063 189 1067 191
rect 1071 190 1077 194
rect 1063 187 1064 189
rect 1066 187 1067 189
rect 1063 186 1067 187
rect 1063 182 1070 186
rect 1013 177 1019 179
rect 1013 175 1014 177
rect 1016 175 1019 177
rect 1013 173 1019 175
rect 1023 177 1027 182
rect 1023 175 1024 177
rect 1026 175 1027 177
rect 1023 173 1027 175
rect 1015 170 1019 173
rect 1015 166 1035 170
rect 1031 162 1035 166
rect 1066 171 1070 182
rect 1073 180 1077 190
rect 1073 178 1074 180
rect 1076 178 1077 180
rect 1073 176 1077 178
rect 1066 170 1084 171
rect 1046 168 1050 170
rect 1066 169 1080 170
rect 1046 166 1047 168
rect 1049 166 1050 168
rect 1031 161 1041 162
rect 1031 159 1037 161
rect 1039 159 1041 161
rect 1031 158 1041 159
rect 1046 161 1050 166
rect 1055 168 1080 169
rect 1082 168 1084 170
rect 1055 166 1057 168
rect 1059 167 1084 168
rect 1059 166 1070 167
rect 1055 165 1070 166
rect 1109 194 1113 198
rect 1109 190 1124 194
rect 1099 181 1105 182
rect 1120 177 1124 190
rect 1127 187 1128 198
rect 1120 175 1121 177
rect 1123 175 1124 177
rect 1120 169 1124 175
rect 1106 168 1124 169
rect 1106 166 1108 168
rect 1110 166 1124 168
rect 1106 165 1124 166
rect 1046 159 1047 161
rect 1049 160 1071 161
rect 1049 159 1067 160
rect 1046 158 1067 159
rect 1069 158 1071 160
rect 937 157 962 158
rect 1046 157 1071 158
rect 1076 157 1080 159
rect -204 155 -203 157
rect -201 155 -200 157
rect -56 155 -55 157
rect -53 155 -52 157
rect -204 152 -200 155
rect -148 154 -142 155
rect -148 152 -146 154
rect -144 152 -142 154
rect -114 154 -108 155
rect -114 152 -112 154
rect -110 152 -108 154
rect -56 152 -52 155
rect -36 155 -30 156
rect -36 153 -34 155
rect -32 153 -30 155
rect -36 152 -30 153
rect -17 155 -11 156
rect -17 153 -15 155
rect -13 153 -11 155
rect -17 152 -11 153
rect 98 155 99 157
rect 101 155 102 157
rect 246 155 247 157
rect 249 155 250 157
rect 98 152 102 155
rect 154 154 160 155
rect 154 152 156 154
rect 158 152 160 154
rect 188 154 194 155
rect 188 152 190 154
rect 192 152 194 154
rect 246 152 250 155
rect 266 155 272 156
rect 266 153 268 155
rect 270 153 272 155
rect 266 152 272 153
rect 285 155 291 156
rect 285 153 287 155
rect 289 153 291 155
rect 285 152 291 153
rect 375 155 376 157
rect 378 155 379 157
rect 523 155 524 157
rect 526 155 527 157
rect 375 152 379 155
rect 431 154 437 155
rect 431 152 433 154
rect 435 152 437 154
rect 465 154 471 155
rect 465 152 467 154
rect 469 152 471 154
rect 523 152 527 155
rect 543 155 549 156
rect 543 153 545 155
rect 547 153 549 155
rect 543 152 549 153
rect 562 155 568 156
rect 562 153 564 155
rect 566 153 568 155
rect 562 152 568 153
rect 651 155 652 157
rect 654 155 655 157
rect 799 155 800 157
rect 802 155 803 157
rect 651 152 655 155
rect 707 154 713 155
rect 707 152 709 154
rect 711 152 713 154
rect 741 154 747 155
rect 741 152 743 154
rect 745 152 747 154
rect 799 152 803 155
rect 819 155 825 156
rect 819 153 821 155
rect 823 153 825 155
rect 819 152 825 153
rect 838 155 844 156
rect 838 153 840 155
rect 842 153 844 155
rect 838 152 844 153
rect 928 155 929 157
rect 931 155 932 157
rect 1076 155 1077 157
rect 1079 155 1080 157
rect 928 152 932 155
rect 984 154 990 155
rect 984 152 986 154
rect 988 152 990 154
rect 1018 154 1024 155
rect 1018 152 1020 154
rect 1022 152 1024 154
rect 1076 152 1080 155
rect 1096 155 1102 156
rect 1096 153 1098 155
rect 1100 153 1102 155
rect 1096 152 1102 153
rect 1115 155 1121 156
rect 1115 153 1117 155
rect 1119 153 1121 155
rect 1115 152 1121 153
rect -269 130 -263 136
rect -204 133 -200 136
rect -148 134 -146 136
rect -144 134 -142 136
rect -148 133 -142 134
rect -114 134 -112 136
rect -110 134 -108 136
rect -114 133 -108 134
rect -56 133 -52 136
rect -204 131 -203 133
rect -201 131 -200 133
rect -56 131 -55 133
rect -53 131 -52 133
rect -36 135 -30 136
rect -36 133 -34 135
rect -32 133 -30 135
rect -36 132 -30 133
rect -17 135 -11 136
rect -17 133 -15 135
rect -13 133 -11 135
rect -17 132 -11 133
rect 98 133 102 136
rect 154 134 156 136
rect 158 134 160 136
rect 154 133 160 134
rect 188 134 190 136
rect 192 134 194 136
rect 188 133 194 134
rect 246 133 250 136
rect 98 131 99 133
rect 101 131 102 133
rect 246 131 247 133
rect 249 131 250 133
rect 266 135 272 136
rect 266 133 268 135
rect 270 133 272 135
rect 266 132 272 133
rect 285 135 291 136
rect 285 133 287 135
rect 289 133 291 135
rect 285 132 291 133
rect 375 133 379 136
rect 431 134 433 136
rect 435 134 437 136
rect 431 133 437 134
rect 465 134 467 136
rect 469 134 471 136
rect 465 133 471 134
rect 523 133 527 136
rect 375 131 376 133
rect 378 131 379 133
rect 523 131 524 133
rect 526 131 527 133
rect 543 135 549 136
rect 543 133 545 135
rect 547 133 549 135
rect 543 132 549 133
rect 562 135 568 136
rect 562 133 564 135
rect 566 133 568 135
rect 562 132 568 133
rect 651 133 655 136
rect 707 134 709 136
rect 711 134 713 136
rect 707 133 713 134
rect 741 134 743 136
rect 745 134 747 136
rect 741 133 747 134
rect 799 133 803 136
rect 651 131 652 133
rect 654 131 655 133
rect 799 131 800 133
rect 802 131 803 133
rect 819 135 825 136
rect 819 133 821 135
rect 823 133 825 135
rect 819 132 825 133
rect 838 135 844 136
rect 838 133 840 135
rect 842 133 844 135
rect 838 132 844 133
rect 928 133 932 136
rect 984 134 986 136
rect 988 134 990 136
rect 984 133 990 134
rect 1018 134 1020 136
rect 1022 134 1024 136
rect 1018 133 1024 134
rect 1076 133 1080 136
rect 928 131 929 133
rect 931 131 932 133
rect 1076 131 1077 133
rect 1079 131 1080 133
rect 1096 135 1102 136
rect 1096 133 1098 135
rect 1100 133 1102 135
rect 1096 132 1102 133
rect 1115 135 1121 136
rect 1115 133 1117 135
rect 1119 133 1121 135
rect 1115 132 1121 133
rect -269 128 -267 130
rect -265 128 -263 130
rect -269 127 -263 128
rect -256 127 -252 129
rect -256 125 -255 127
rect -253 125 -252 127
rect -282 122 -278 124
rect -282 120 -281 122
rect -279 120 -278 122
rect -282 114 -278 120
rect -256 122 -252 125
rect -256 118 -232 122
rect -282 110 -271 114
rect -275 104 -271 110
rect -236 114 -232 118
rect -256 113 -240 114
rect -256 111 -244 113
rect -242 111 -240 113
rect -256 110 -240 111
rect -236 112 -231 114
rect -236 110 -234 112
rect -232 110 -231 112
rect -256 104 -252 110
rect -236 108 -231 110
rect -236 106 -232 108
rect -275 103 -252 104
rect -275 101 -273 103
rect -271 101 -252 103
rect -275 100 -252 101
rect -264 89 -260 91
rect -264 87 -263 89
rect -261 87 -260 89
rect -264 82 -260 87
rect -256 89 -252 100
rect -248 103 -232 106
rect -248 101 -247 103
rect -245 102 -232 103
rect -245 101 -244 102
rect -248 96 -244 101
rect -248 94 -247 96
rect -245 94 -244 96
rect -248 92 -244 94
rect -204 129 -200 131
rect -195 130 -170 131
rect -86 130 -61 131
rect -195 128 -193 130
rect -191 129 -170 130
rect -191 128 -173 129
rect -195 127 -173 128
rect -171 127 -170 129
rect -194 122 -179 123
rect -194 121 -183 122
rect -208 120 -183 121
rect -181 120 -179 122
rect -208 118 -206 120
rect -204 119 -179 120
rect -174 122 -170 127
rect -165 129 -155 130
rect -165 127 -163 129
rect -161 127 -155 129
rect -165 126 -155 127
rect -174 120 -173 122
rect -171 120 -170 122
rect -204 118 -190 119
rect -174 118 -170 120
rect -208 117 -190 118
rect -201 110 -197 112
rect -201 108 -200 110
rect -198 108 -197 110
rect -201 98 -197 108
rect -194 106 -190 117
rect -159 122 -155 126
rect -159 118 -139 122
rect -143 115 -139 118
rect -151 113 -147 115
rect -151 111 -150 113
rect -148 111 -147 113
rect -151 106 -147 111
rect -143 113 -137 115
rect -143 111 -140 113
rect -138 111 -137 113
rect -143 109 -137 111
rect -194 102 -187 106
rect -191 101 -187 102
rect -191 99 -190 101
rect -188 99 -187 101
rect -201 94 -195 98
rect -191 97 -187 99
rect -143 98 -139 109
rect -179 97 -139 98
rect -179 95 -155 97
rect -153 95 -139 97
rect -179 94 -139 95
rect -199 90 -175 94
rect -156 90 -152 94
rect -101 129 -91 130
rect -101 127 -95 129
rect -93 127 -91 129
rect -101 126 -91 127
rect -86 129 -65 130
rect -86 127 -85 129
rect -83 128 -65 129
rect -63 128 -61 130
rect -56 129 -52 131
rect -83 127 -61 128
rect -101 122 -97 126
rect -117 118 -97 122
rect -117 115 -113 118
rect -119 113 -113 115
rect -119 111 -118 113
rect -116 111 -113 113
rect -119 109 -113 111
rect -117 98 -113 109
rect -109 113 -105 115
rect -86 122 -82 127
rect 7 129 27 130
rect 7 127 9 129
rect 11 127 27 129
rect 7 126 27 127
rect -86 120 -85 122
rect -83 120 -82 122
rect -86 118 -82 120
rect -77 122 -62 123
rect -77 120 -75 122
rect -73 121 -62 122
rect -73 120 -48 121
rect -77 119 -52 120
rect -66 118 -52 119
rect -50 118 -48 120
rect -66 117 -48 118
rect -109 111 -108 113
rect -106 111 -105 113
rect -109 106 -105 111
rect -66 106 -62 117
rect -69 102 -62 106
rect -59 110 -55 112
rect -59 108 -58 110
rect -56 108 -55 110
rect -69 101 -65 102
rect -69 99 -68 101
rect -66 99 -65 101
rect -117 97 -77 98
rect -69 97 -65 99
rect -59 98 -55 108
rect -26 122 -8 123
rect -26 120 -24 122
rect -22 120 -8 122
rect -26 119 -8 120
rect -12 113 -8 119
rect -12 111 -11 113
rect -9 111 -8 113
rect -33 106 -27 107
rect -117 95 -103 97
rect -101 95 -77 97
rect -117 94 -77 95
rect -61 94 -55 98
rect -104 90 -100 94
rect -81 90 -57 94
rect -12 98 -8 111
rect 23 122 27 126
rect 47 129 67 130
rect 47 127 49 129
rect 51 127 67 129
rect 47 126 67 127
rect 38 123 39 125
rect 23 118 35 122
rect 31 113 35 118
rect 31 111 32 113
rect 34 111 35 113
rect -23 94 -8 98
rect -23 90 -19 94
rect -5 90 -4 101
rect 31 99 35 111
rect 63 122 67 126
rect 78 123 79 125
rect 63 118 75 122
rect 71 113 75 118
rect 71 111 72 113
rect 74 111 75 113
rect 18 96 35 99
rect 18 94 19 96
rect 21 95 35 96
rect 21 94 22 95
rect -169 89 -163 90
rect -256 88 -223 89
rect -256 86 -227 88
rect -225 86 -223 88
rect -256 85 -223 86
rect -169 87 -167 89
rect -165 87 -163 89
rect -264 80 -263 82
rect -261 80 -260 82
rect -204 82 -198 83
rect -204 80 -202 82
rect -200 80 -198 82
rect -169 82 -163 87
rect -156 88 -155 90
rect -153 88 -152 90
rect -156 86 -152 88
rect -147 89 -141 90
rect -147 87 -145 89
rect -143 87 -141 89
rect -169 80 -167 82
rect -165 80 -163 82
rect -147 82 -141 87
rect -147 80 -145 82
rect -143 80 -141 82
rect -115 89 -109 90
rect -115 87 -113 89
rect -111 87 -109 89
rect -115 82 -109 87
rect -104 88 -103 90
rect -101 88 -100 90
rect -104 86 -100 88
rect -93 89 -87 90
rect -93 87 -91 89
rect -89 87 -87 89
rect -115 80 -113 82
rect -111 80 -109 82
rect -93 82 -87 87
rect -36 89 -19 90
rect -36 87 -34 89
rect -32 87 -19 89
rect -36 86 -19 87
rect 7 89 13 90
rect 7 87 9 89
rect 11 87 13 89
rect -93 80 -91 82
rect -89 80 -87 82
rect -58 82 -52 83
rect -58 80 -56 82
rect -54 80 -52 82
rect -17 82 -11 83
rect -17 80 -15 82
rect -13 80 -11 82
rect 7 80 13 87
rect 18 89 22 94
rect 71 99 75 111
rect 58 96 75 99
rect 58 94 59 96
rect 61 95 75 96
rect 61 94 62 95
rect 18 87 19 89
rect 21 87 22 89
rect 18 85 22 87
rect 27 91 33 92
rect 27 89 29 91
rect 31 89 33 91
rect 47 89 53 90
rect 27 80 33 89
rect 47 87 49 89
rect 51 87 53 89
rect 47 80 53 87
rect 58 89 62 94
rect 98 129 102 131
rect 107 130 132 131
rect 216 130 241 131
rect 107 128 109 130
rect 111 129 132 130
rect 111 128 129 129
rect 107 127 129 128
rect 131 127 132 129
rect 108 122 123 123
rect 108 121 119 122
rect 94 120 119 121
rect 121 120 123 122
rect 94 118 96 120
rect 98 119 123 120
rect 128 122 132 127
rect 137 129 147 130
rect 137 127 139 129
rect 141 127 147 129
rect 137 126 147 127
rect 128 120 129 122
rect 131 120 132 122
rect 98 118 112 119
rect 128 118 132 120
rect 94 117 112 118
rect 101 110 105 112
rect 101 108 102 110
rect 104 108 105 110
rect 101 98 105 108
rect 108 106 112 117
rect 143 122 147 126
rect 143 118 163 122
rect 159 115 163 118
rect 151 113 155 115
rect 151 111 152 113
rect 154 111 155 113
rect 151 106 155 111
rect 159 113 165 115
rect 159 111 162 113
rect 164 111 165 113
rect 159 109 165 111
rect 108 102 115 106
rect 111 101 115 102
rect 111 99 112 101
rect 114 99 115 101
rect 101 94 107 98
rect 111 97 115 99
rect 159 98 163 109
rect 123 97 163 98
rect 123 95 147 97
rect 149 95 163 97
rect 123 94 163 95
rect 58 87 59 89
rect 61 87 62 89
rect 58 85 62 87
rect 67 91 73 92
rect 67 89 69 91
rect 71 89 73 91
rect 103 90 127 94
rect 146 90 150 94
rect 201 129 211 130
rect 201 127 207 129
rect 209 127 211 129
rect 201 126 211 127
rect 216 129 237 130
rect 216 127 217 129
rect 219 128 237 129
rect 239 128 241 130
rect 246 129 250 131
rect 219 127 241 128
rect 201 122 205 126
rect 185 118 205 122
rect 185 115 189 118
rect 183 113 189 115
rect 183 111 184 113
rect 186 111 189 113
rect 183 109 189 111
rect 185 98 189 109
rect 193 113 197 115
rect 216 122 220 127
rect 314 129 334 130
rect 314 127 316 129
rect 318 127 334 129
rect 314 126 334 127
rect 216 120 217 122
rect 219 120 220 122
rect 216 118 220 120
rect 225 122 240 123
rect 225 120 227 122
rect 229 121 240 122
rect 229 120 254 121
rect 225 119 250 120
rect 236 118 250 119
rect 252 118 254 120
rect 236 117 254 118
rect 193 111 194 113
rect 196 111 197 113
rect 193 106 197 111
rect 236 106 240 117
rect 233 102 240 106
rect 243 110 247 112
rect 243 108 244 110
rect 246 108 247 110
rect 233 101 237 102
rect 233 99 234 101
rect 236 99 237 101
rect 185 97 225 98
rect 233 97 237 99
rect 243 98 247 108
rect 276 122 294 123
rect 276 120 278 122
rect 280 120 294 122
rect 276 119 294 120
rect 290 113 294 119
rect 290 111 291 113
rect 293 111 294 113
rect 269 106 275 107
rect 185 95 199 97
rect 201 95 225 97
rect 185 94 225 95
rect 241 94 247 98
rect 198 90 202 94
rect 221 90 245 94
rect 290 98 294 111
rect 279 94 294 98
rect 279 90 283 94
rect 297 90 298 101
rect 330 122 334 126
rect 345 123 346 125
rect 330 118 342 122
rect 338 113 342 118
rect 338 111 339 113
rect 341 111 342 113
rect 338 99 342 111
rect 325 96 342 99
rect 325 94 326 96
rect 328 95 342 96
rect 328 94 329 95
rect 67 80 73 89
rect 133 89 139 90
rect 133 87 135 89
rect 137 87 139 89
rect 98 82 104 83
rect 98 80 100 82
rect 102 80 104 82
rect 133 82 139 87
rect 146 88 147 90
rect 149 88 150 90
rect 146 86 150 88
rect 155 89 161 90
rect 155 87 157 89
rect 159 87 161 89
rect 133 80 135 82
rect 137 80 139 82
rect 155 82 161 87
rect 155 80 157 82
rect 159 80 161 82
rect 187 89 193 90
rect 187 87 189 89
rect 191 87 193 89
rect 187 82 193 87
rect 198 88 199 90
rect 201 88 202 90
rect 198 86 202 88
rect 209 89 215 90
rect 209 87 211 89
rect 213 87 215 89
rect 187 80 189 82
rect 191 80 193 82
rect 209 82 215 87
rect 266 89 283 90
rect 266 87 268 89
rect 270 87 283 89
rect 266 86 283 87
rect 314 89 320 90
rect 314 87 316 89
rect 318 87 320 89
rect 209 80 211 82
rect 213 80 215 82
rect 244 82 250 83
rect 244 80 246 82
rect 248 80 250 82
rect 285 82 291 83
rect 285 80 287 82
rect 289 80 291 82
rect 314 80 320 87
rect 325 89 329 94
rect 375 129 379 131
rect 384 130 409 131
rect 493 130 518 131
rect 384 128 386 130
rect 388 129 409 130
rect 388 128 406 129
rect 384 127 406 128
rect 408 127 409 129
rect 385 122 400 123
rect 385 121 396 122
rect 371 120 396 121
rect 398 120 400 122
rect 371 118 373 120
rect 375 119 400 120
rect 405 122 409 127
rect 414 129 424 130
rect 414 127 416 129
rect 418 127 424 129
rect 414 126 424 127
rect 405 120 406 122
rect 408 120 409 122
rect 375 118 389 119
rect 405 118 409 120
rect 371 117 389 118
rect 378 110 382 112
rect 378 108 379 110
rect 381 108 382 110
rect 378 98 382 108
rect 385 106 389 117
rect 420 122 424 126
rect 420 118 440 122
rect 436 115 440 118
rect 428 113 432 115
rect 428 111 429 113
rect 431 111 432 113
rect 428 106 432 111
rect 436 113 442 115
rect 436 111 439 113
rect 441 111 442 113
rect 436 109 442 111
rect 385 102 392 106
rect 388 101 392 102
rect 388 99 389 101
rect 391 99 392 101
rect 378 94 384 98
rect 388 97 392 99
rect 436 98 440 109
rect 400 97 440 98
rect 400 95 424 97
rect 426 95 440 97
rect 400 94 440 95
rect 325 87 326 89
rect 328 87 329 89
rect 325 85 329 87
rect 334 91 340 92
rect 334 89 336 91
rect 338 89 340 91
rect 380 90 404 94
rect 423 90 427 94
rect 478 129 488 130
rect 478 127 484 129
rect 486 127 488 129
rect 478 126 488 127
rect 493 129 514 130
rect 493 127 494 129
rect 496 128 514 129
rect 516 128 518 130
rect 523 129 527 131
rect 496 127 518 128
rect 478 122 482 126
rect 462 118 482 122
rect 462 115 466 118
rect 460 113 466 115
rect 460 111 461 113
rect 463 111 466 113
rect 460 109 466 111
rect 462 98 466 109
rect 470 113 474 115
rect 493 122 497 127
rect 591 129 611 130
rect 591 127 593 129
rect 595 127 611 129
rect 591 126 611 127
rect 493 120 494 122
rect 496 120 497 122
rect 493 118 497 120
rect 502 122 517 123
rect 502 120 504 122
rect 506 121 517 122
rect 506 120 531 121
rect 502 119 527 120
rect 513 118 527 119
rect 529 118 531 120
rect 513 117 531 118
rect 470 111 471 113
rect 473 111 474 113
rect 470 106 474 111
rect 513 106 517 117
rect 510 102 517 106
rect 520 110 524 112
rect 520 108 521 110
rect 523 108 524 110
rect 510 101 514 102
rect 510 99 511 101
rect 513 99 514 101
rect 462 97 502 98
rect 510 97 514 99
rect 520 98 524 108
rect 553 122 571 123
rect 553 120 555 122
rect 557 120 571 122
rect 553 119 571 120
rect 567 113 571 119
rect 567 111 568 113
rect 570 111 571 113
rect 546 106 552 107
rect 462 95 476 97
rect 478 95 502 97
rect 462 94 502 95
rect 518 94 524 98
rect 475 90 479 94
rect 498 90 522 94
rect 567 98 571 111
rect 556 94 571 98
rect 556 90 560 94
rect 574 90 575 101
rect 607 122 611 126
rect 622 123 623 125
rect 607 118 619 122
rect 615 113 619 118
rect 615 111 616 113
rect 618 111 619 113
rect 615 99 619 111
rect 602 96 619 99
rect 602 94 603 96
rect 605 95 619 96
rect 605 94 606 95
rect 334 80 340 89
rect 410 89 416 90
rect 410 87 412 89
rect 414 87 416 89
rect 375 82 381 83
rect 375 80 377 82
rect 379 80 381 82
rect 410 82 416 87
rect 423 88 424 90
rect 426 88 427 90
rect 423 86 427 88
rect 432 89 438 90
rect 432 87 434 89
rect 436 87 438 89
rect 410 80 412 82
rect 414 80 416 82
rect 432 82 438 87
rect 432 80 434 82
rect 436 80 438 82
rect 464 89 470 90
rect 464 87 466 89
rect 468 87 470 89
rect 464 82 470 87
rect 475 88 476 90
rect 478 88 479 90
rect 475 86 479 88
rect 486 89 492 90
rect 486 87 488 89
rect 490 87 492 89
rect 464 80 466 82
rect 468 80 470 82
rect 486 82 492 87
rect 543 89 560 90
rect 543 87 545 89
rect 547 87 560 89
rect 543 86 560 87
rect 591 89 597 90
rect 591 87 593 89
rect 595 87 597 89
rect 486 80 488 82
rect 490 80 492 82
rect 521 82 527 83
rect 521 80 523 82
rect 525 80 527 82
rect 562 82 568 83
rect 562 80 564 82
rect 566 80 568 82
rect 591 80 597 87
rect 602 89 606 94
rect 651 129 655 131
rect 660 130 685 131
rect 769 130 794 131
rect 660 128 662 130
rect 664 129 685 130
rect 664 128 682 129
rect 660 127 682 128
rect 684 127 685 129
rect 661 122 676 123
rect 661 121 672 122
rect 647 120 672 121
rect 674 120 676 122
rect 647 118 649 120
rect 651 119 676 120
rect 681 122 685 127
rect 690 129 700 130
rect 690 127 692 129
rect 694 127 700 129
rect 690 126 700 127
rect 681 120 682 122
rect 684 120 685 122
rect 651 118 665 119
rect 681 118 685 120
rect 647 117 665 118
rect 654 110 658 112
rect 654 108 655 110
rect 657 108 658 110
rect 654 98 658 108
rect 661 106 665 117
rect 696 122 700 126
rect 696 118 716 122
rect 712 115 716 118
rect 704 113 708 115
rect 704 111 705 113
rect 707 111 708 113
rect 704 106 708 111
rect 712 113 718 115
rect 712 111 715 113
rect 717 111 718 113
rect 712 109 718 111
rect 661 102 668 106
rect 664 101 668 102
rect 664 99 665 101
rect 667 99 668 101
rect 654 94 660 98
rect 664 97 668 99
rect 712 98 716 109
rect 676 97 716 98
rect 676 95 700 97
rect 702 95 716 97
rect 676 94 716 95
rect 602 87 603 89
rect 605 87 606 89
rect 602 85 606 87
rect 611 91 617 92
rect 611 89 613 91
rect 615 89 617 91
rect 656 90 680 94
rect 699 90 703 94
rect 754 129 764 130
rect 754 127 760 129
rect 762 127 764 129
rect 754 126 764 127
rect 769 129 790 130
rect 769 127 770 129
rect 772 128 790 129
rect 792 128 794 130
rect 799 129 803 131
rect 772 127 794 128
rect 754 122 758 126
rect 738 118 758 122
rect 738 115 742 118
rect 736 113 742 115
rect 736 111 737 113
rect 739 111 742 113
rect 736 109 742 111
rect 738 98 742 109
rect 746 113 750 115
rect 769 122 773 127
rect 867 129 887 130
rect 867 127 869 129
rect 871 127 887 129
rect 867 126 887 127
rect 769 120 770 122
rect 772 120 773 122
rect 769 118 773 120
rect 778 122 793 123
rect 778 120 780 122
rect 782 121 793 122
rect 782 120 807 121
rect 778 119 803 120
rect 789 118 803 119
rect 805 118 807 120
rect 789 117 807 118
rect 746 111 747 113
rect 749 111 750 113
rect 746 106 750 111
rect 789 106 793 117
rect 786 102 793 106
rect 796 110 800 112
rect 796 108 797 110
rect 799 108 800 110
rect 786 101 790 102
rect 786 99 787 101
rect 789 99 790 101
rect 738 97 778 98
rect 786 97 790 99
rect 796 98 800 108
rect 829 122 847 123
rect 829 120 831 122
rect 833 120 847 122
rect 829 119 847 120
rect 843 113 847 119
rect 843 111 844 113
rect 846 111 847 113
rect 822 106 828 107
rect 738 95 752 97
rect 754 95 778 97
rect 738 94 778 95
rect 794 94 800 98
rect 751 90 755 94
rect 774 90 798 94
rect 843 98 847 111
rect 832 94 847 98
rect 832 90 836 94
rect 850 90 851 101
rect 883 122 887 126
rect 898 123 899 125
rect 883 118 895 122
rect 891 113 895 118
rect 891 111 892 113
rect 894 111 895 113
rect 891 99 895 111
rect 878 96 895 99
rect 878 94 879 96
rect 881 95 895 96
rect 881 94 882 95
rect 611 80 617 89
rect 686 89 692 90
rect 686 87 688 89
rect 690 87 692 89
rect 651 82 657 83
rect 651 80 653 82
rect 655 80 657 82
rect 686 82 692 87
rect 699 88 700 90
rect 702 88 703 90
rect 699 86 703 88
rect 708 89 714 90
rect 708 87 710 89
rect 712 87 714 89
rect 686 80 688 82
rect 690 80 692 82
rect 708 82 714 87
rect 708 80 710 82
rect 712 80 714 82
rect 740 89 746 90
rect 740 87 742 89
rect 744 87 746 89
rect 740 82 746 87
rect 751 88 752 90
rect 754 88 755 90
rect 751 86 755 88
rect 762 89 768 90
rect 762 87 764 89
rect 766 87 768 89
rect 740 80 742 82
rect 744 80 746 82
rect 762 82 768 87
rect 819 89 836 90
rect 819 87 821 89
rect 823 87 836 89
rect 819 86 836 87
rect 867 89 873 90
rect 867 87 869 89
rect 871 87 873 89
rect 762 80 764 82
rect 766 80 768 82
rect 797 82 803 83
rect 797 80 799 82
rect 801 80 803 82
rect 838 82 844 83
rect 838 80 840 82
rect 842 80 844 82
rect 867 80 873 87
rect 878 89 882 94
rect 928 129 932 131
rect 937 130 962 131
rect 1046 130 1071 131
rect 937 128 939 130
rect 941 129 962 130
rect 941 128 959 129
rect 937 127 959 128
rect 961 127 962 129
rect 938 122 953 123
rect 938 121 949 122
rect 924 120 949 121
rect 951 120 953 122
rect 924 118 926 120
rect 928 119 953 120
rect 958 122 962 127
rect 967 129 977 130
rect 967 127 969 129
rect 971 127 977 129
rect 967 126 977 127
rect 958 120 959 122
rect 961 120 962 122
rect 928 118 942 119
rect 958 118 962 120
rect 924 117 942 118
rect 931 110 935 112
rect 931 108 932 110
rect 934 108 935 110
rect 931 98 935 108
rect 938 106 942 117
rect 973 122 977 126
rect 973 118 993 122
rect 989 115 993 118
rect 981 113 985 115
rect 981 111 982 113
rect 984 111 985 113
rect 981 106 985 111
rect 989 113 995 115
rect 989 111 992 113
rect 994 111 995 113
rect 989 109 995 111
rect 938 102 945 106
rect 941 101 945 102
rect 941 99 942 101
rect 944 99 945 101
rect 931 94 937 98
rect 941 97 945 99
rect 989 98 993 109
rect 953 97 993 98
rect 953 95 977 97
rect 979 95 993 97
rect 953 94 993 95
rect 878 87 879 89
rect 881 87 882 89
rect 878 85 882 87
rect 887 91 893 92
rect 887 89 889 91
rect 891 89 893 91
rect 933 90 957 94
rect 976 90 980 94
rect 1031 129 1041 130
rect 1031 127 1037 129
rect 1039 127 1041 129
rect 1031 126 1041 127
rect 1046 129 1067 130
rect 1046 127 1047 129
rect 1049 128 1067 129
rect 1069 128 1071 130
rect 1076 129 1080 131
rect 1049 127 1071 128
rect 1031 122 1035 126
rect 1015 118 1035 122
rect 1015 115 1019 118
rect 1013 113 1019 115
rect 1013 111 1014 113
rect 1016 111 1019 113
rect 1013 109 1019 111
rect 1015 98 1019 109
rect 1023 113 1027 115
rect 1046 122 1050 127
rect 1046 120 1047 122
rect 1049 120 1050 122
rect 1046 118 1050 120
rect 1055 122 1070 123
rect 1055 120 1057 122
rect 1059 121 1070 122
rect 1059 120 1084 121
rect 1055 119 1080 120
rect 1066 118 1080 119
rect 1082 118 1084 120
rect 1066 117 1084 118
rect 1023 111 1024 113
rect 1026 111 1027 113
rect 1023 106 1027 111
rect 1066 106 1070 117
rect 1063 102 1070 106
rect 1073 110 1077 112
rect 1073 108 1074 110
rect 1076 108 1077 110
rect 1063 101 1067 102
rect 1063 99 1064 101
rect 1066 99 1067 101
rect 1015 97 1055 98
rect 1063 97 1067 99
rect 1073 98 1077 108
rect 1106 122 1124 123
rect 1106 120 1108 122
rect 1110 120 1124 122
rect 1106 119 1124 120
rect 1120 113 1124 119
rect 1120 111 1121 113
rect 1123 111 1124 113
rect 1099 106 1105 107
rect 1015 95 1029 97
rect 1031 95 1055 97
rect 1015 94 1055 95
rect 1071 94 1077 98
rect 1028 90 1032 94
rect 1051 90 1075 94
rect 1120 98 1124 111
rect 1109 94 1124 98
rect 1109 90 1113 94
rect 1127 90 1128 101
rect 887 80 893 89
rect 963 89 969 90
rect 963 87 965 89
rect 967 87 969 89
rect 928 82 934 83
rect 928 80 930 82
rect 932 80 934 82
rect 963 82 969 87
rect 976 88 977 90
rect 979 88 980 90
rect 976 86 980 88
rect 985 89 991 90
rect 985 87 987 89
rect 989 87 991 89
rect 963 80 965 82
rect 967 80 969 82
rect 985 82 991 87
rect 985 80 987 82
rect 989 80 991 82
rect 1017 89 1023 90
rect 1017 87 1019 89
rect 1021 87 1023 89
rect 1017 82 1023 87
rect 1028 88 1029 90
rect 1031 88 1032 90
rect 1028 86 1032 88
rect 1039 89 1045 90
rect 1039 87 1041 89
rect 1043 87 1045 89
rect 1017 80 1019 82
rect 1021 80 1023 82
rect 1039 82 1045 87
rect 1096 89 1113 90
rect 1096 87 1098 89
rect 1100 87 1113 89
rect 1096 86 1113 87
rect 1039 80 1041 82
rect 1043 80 1045 82
rect 1074 82 1080 83
rect 1074 80 1076 82
rect 1078 80 1080 82
rect 1115 82 1121 83
rect 1115 80 1117 82
rect 1119 80 1121 82
rect -264 62 -263 64
rect -261 62 -260 64
rect -264 57 -260 62
rect -204 62 -202 64
rect -200 62 -198 64
rect -204 61 -198 62
rect -169 62 -167 64
rect -165 62 -163 64
rect -264 55 -263 57
rect -261 55 -260 57
rect -264 53 -260 55
rect -256 58 -223 59
rect -256 56 -227 58
rect -225 56 -223 58
rect -256 55 -223 56
rect -169 57 -163 62
rect -147 62 -145 64
rect -143 62 -141 64
rect -169 55 -167 57
rect -165 55 -163 57
rect -256 44 -252 55
rect -169 54 -163 55
rect -156 56 -152 58
rect -156 54 -155 56
rect -153 54 -152 56
rect -147 57 -141 62
rect -147 55 -145 57
rect -143 55 -141 57
rect -147 54 -141 55
rect -115 62 -113 64
rect -111 62 -109 64
rect -115 57 -109 62
rect -93 62 -91 64
rect -89 62 -87 64
rect -115 55 -113 57
rect -111 55 -109 57
rect -115 54 -109 55
rect -104 56 -100 58
rect -104 54 -103 56
rect -101 54 -100 56
rect -93 57 -87 62
rect -58 62 -56 64
rect -54 62 -52 64
rect -58 61 -52 62
rect -17 62 -15 64
rect -13 62 -11 64
rect -17 61 -11 62
rect -93 55 -91 57
rect -89 55 -87 57
rect -93 54 -87 55
rect -36 57 -19 58
rect -36 55 -34 57
rect -32 55 -19 57
rect -36 54 -19 55
rect 7 57 13 64
rect 7 55 9 57
rect 11 55 13 57
rect 7 54 13 55
rect 18 57 22 59
rect 18 55 19 57
rect 21 55 22 57
rect -275 43 -252 44
rect -275 41 -273 43
rect -271 41 -252 43
rect -275 40 -252 41
rect -275 34 -271 40
rect -282 30 -271 34
rect -282 24 -278 30
rect -256 34 -252 40
rect -248 50 -244 52
rect -248 48 -247 50
rect -245 48 -244 50
rect -248 43 -244 48
rect -248 41 -247 43
rect -245 42 -244 43
rect -245 41 -232 42
rect -248 38 -232 41
rect -236 36 -232 38
rect -236 34 -231 36
rect -256 33 -240 34
rect -256 31 -244 33
rect -242 31 -240 33
rect -256 30 -240 31
rect -236 32 -234 34
rect -232 32 -231 34
rect -236 30 -231 32
rect -282 22 -281 24
rect -279 22 -278 24
rect -282 20 -278 22
rect -236 26 -232 30
rect -256 22 -232 26
rect -256 19 -252 22
rect -256 17 -255 19
rect -253 17 -252 19
rect -269 16 -263 17
rect -269 14 -267 16
rect -265 14 -263 16
rect -256 15 -252 17
rect -199 50 -175 54
rect -156 50 -152 54
rect -201 46 -195 50
rect -179 49 -139 50
rect -179 47 -155 49
rect -153 47 -139 49
rect -201 36 -197 46
rect -191 45 -187 47
rect -179 46 -139 47
rect -191 43 -190 45
rect -188 43 -187 45
rect -191 42 -187 43
rect -201 34 -200 36
rect -198 34 -197 36
rect -201 32 -197 34
rect -194 38 -187 42
rect -194 27 -190 38
rect -151 33 -147 38
rect -151 31 -150 33
rect -148 31 -147 33
rect -208 26 -190 27
rect -208 24 -206 26
rect -204 25 -190 26
rect -204 24 -179 25
rect -208 23 -183 24
rect -194 22 -183 23
rect -181 22 -179 24
rect -194 21 -179 22
rect -174 24 -170 26
rect -174 22 -173 24
rect -171 22 -170 24
rect -174 17 -170 22
rect -151 29 -147 31
rect -143 35 -139 46
rect -143 33 -137 35
rect -143 31 -140 33
rect -138 31 -137 33
rect -143 29 -137 31
rect -143 26 -139 29
rect -159 22 -139 26
rect -159 18 -155 22
rect -195 16 -173 17
rect -269 8 -263 14
rect -204 13 -200 15
rect -195 14 -193 16
rect -191 15 -173 16
rect -171 15 -170 17
rect -191 14 -170 15
rect -165 17 -155 18
rect -165 15 -163 17
rect -161 15 -155 17
rect -165 14 -155 15
rect -104 50 -100 54
rect -81 50 -57 54
rect -117 49 -77 50
rect -117 47 -103 49
rect -101 47 -77 49
rect -117 46 -77 47
rect -117 35 -113 46
rect -69 45 -65 47
rect -61 46 -55 50
rect -69 43 -68 45
rect -66 43 -65 45
rect -69 42 -65 43
rect -69 38 -62 42
rect -119 33 -113 35
rect -119 31 -118 33
rect -116 31 -113 33
rect -119 29 -113 31
rect -109 33 -105 38
rect -109 31 -108 33
rect -106 31 -105 33
rect -109 29 -105 31
rect -117 26 -113 29
rect -117 22 -97 26
rect -101 18 -97 22
rect -66 27 -62 38
rect -59 36 -55 46
rect -59 34 -58 36
rect -56 34 -55 36
rect -59 32 -55 34
rect -66 26 -48 27
rect -86 24 -82 26
rect -66 25 -52 26
rect -86 22 -85 24
rect -83 22 -82 24
rect -101 17 -91 18
rect -101 15 -95 17
rect -93 15 -91 17
rect -101 14 -91 15
rect -86 17 -82 22
rect -77 24 -52 25
rect -50 24 -48 26
rect -77 22 -75 24
rect -73 23 -48 24
rect -73 22 -62 23
rect -77 21 -62 22
rect -23 50 -19 54
rect -23 46 -8 50
rect -33 37 -27 38
rect -12 33 -8 46
rect -5 43 -4 54
rect -12 31 -11 33
rect -9 31 -8 33
rect -12 25 -8 31
rect 18 50 22 55
rect 27 55 33 64
rect 27 53 29 55
rect 31 53 33 55
rect 47 57 53 64
rect 47 55 49 57
rect 51 55 53 57
rect 47 54 53 55
rect 58 57 62 59
rect 58 55 59 57
rect 61 55 62 57
rect 27 52 33 53
rect 18 48 19 50
rect 21 49 22 50
rect 21 48 35 49
rect 18 45 35 48
rect -26 24 -8 25
rect -26 22 -24 24
rect -22 22 -8 24
rect -26 21 -8 22
rect 31 33 35 45
rect 31 31 32 33
rect 34 31 35 33
rect 31 26 35 31
rect 23 22 35 26
rect 23 18 27 22
rect 38 19 39 21
rect 58 50 62 55
rect 67 55 73 64
rect 98 62 100 64
rect 102 62 104 64
rect 98 61 104 62
rect 133 62 135 64
rect 137 62 139 64
rect 67 53 69 55
rect 71 53 73 55
rect 133 57 139 62
rect 155 62 157 64
rect 159 62 161 64
rect 133 55 135 57
rect 137 55 139 57
rect 133 54 139 55
rect 146 56 150 58
rect 146 54 147 56
rect 149 54 150 56
rect 155 57 161 62
rect 155 55 157 57
rect 159 55 161 57
rect 155 54 161 55
rect 187 62 189 64
rect 191 62 193 64
rect 187 57 193 62
rect 209 62 211 64
rect 213 62 215 64
rect 187 55 189 57
rect 191 55 193 57
rect 187 54 193 55
rect 198 56 202 58
rect 198 54 199 56
rect 201 54 202 56
rect 209 57 215 62
rect 244 62 246 64
rect 248 62 250 64
rect 244 61 250 62
rect 285 62 287 64
rect 289 62 291 64
rect 285 61 291 62
rect 209 55 211 57
rect 213 55 215 57
rect 209 54 215 55
rect 266 57 283 58
rect 266 55 268 57
rect 270 55 283 57
rect 266 54 283 55
rect 314 57 320 64
rect 314 55 316 57
rect 318 55 320 57
rect 314 54 320 55
rect 325 57 329 59
rect 325 55 326 57
rect 328 55 329 57
rect 67 52 73 53
rect 58 48 59 50
rect 61 49 62 50
rect 61 48 75 49
rect 58 45 75 48
rect 71 33 75 45
rect 71 31 72 33
rect 74 31 75 33
rect 71 26 75 31
rect 63 22 75 26
rect -86 15 -85 17
rect -83 16 -61 17
rect -83 15 -65 16
rect -86 14 -65 15
rect -63 14 -61 16
rect -195 13 -170 14
rect -86 13 -61 14
rect -56 13 -52 15
rect 7 17 27 18
rect 7 15 9 17
rect 11 15 27 17
rect 7 14 27 15
rect 63 18 67 22
rect 78 19 79 21
rect 47 17 67 18
rect 47 15 49 17
rect 51 15 67 17
rect 47 14 67 15
rect 103 50 127 54
rect 146 50 150 54
rect 101 46 107 50
rect 123 49 163 50
rect 123 47 147 49
rect 149 47 163 49
rect 101 36 105 46
rect 111 45 115 47
rect 123 46 163 47
rect 111 43 112 45
rect 114 43 115 45
rect 111 42 115 43
rect 101 34 102 36
rect 104 34 105 36
rect 101 32 105 34
rect 108 38 115 42
rect 108 27 112 38
rect 151 33 155 38
rect 151 31 152 33
rect 154 31 155 33
rect 94 26 112 27
rect 94 24 96 26
rect 98 25 112 26
rect 98 24 123 25
rect 94 23 119 24
rect 108 22 119 23
rect 121 22 123 24
rect 108 21 123 22
rect 128 24 132 26
rect 128 22 129 24
rect 131 22 132 24
rect 128 17 132 22
rect 151 29 155 31
rect 159 35 163 46
rect 159 33 165 35
rect 159 31 162 33
rect 164 31 165 33
rect 159 29 165 31
rect 159 26 163 29
rect 143 22 163 26
rect 143 18 147 22
rect 107 16 129 17
rect 98 13 102 15
rect 107 14 109 16
rect 111 15 129 16
rect 131 15 132 17
rect 111 14 132 15
rect 137 17 147 18
rect 137 15 139 17
rect 141 15 147 17
rect 137 14 147 15
rect 198 50 202 54
rect 221 50 245 54
rect 185 49 225 50
rect 185 47 199 49
rect 201 47 225 49
rect 185 46 225 47
rect 185 35 189 46
rect 233 45 237 47
rect 241 46 247 50
rect 233 43 234 45
rect 236 43 237 45
rect 233 42 237 43
rect 233 38 240 42
rect 183 33 189 35
rect 183 31 184 33
rect 186 31 189 33
rect 183 29 189 31
rect 193 33 197 38
rect 193 31 194 33
rect 196 31 197 33
rect 193 29 197 31
rect 185 26 189 29
rect 185 22 205 26
rect 201 18 205 22
rect 236 27 240 38
rect 243 36 247 46
rect 243 34 244 36
rect 246 34 247 36
rect 243 32 247 34
rect 236 26 254 27
rect 216 24 220 26
rect 236 25 250 26
rect 216 22 217 24
rect 219 22 220 24
rect 201 17 211 18
rect 201 15 207 17
rect 209 15 211 17
rect 201 14 211 15
rect 216 17 220 22
rect 225 24 250 25
rect 252 24 254 26
rect 225 22 227 24
rect 229 23 254 24
rect 279 50 283 54
rect 279 46 294 50
rect 269 37 275 38
rect 229 22 240 23
rect 225 21 240 22
rect 290 33 294 46
rect 297 43 298 54
rect 290 31 291 33
rect 293 31 294 33
rect 290 25 294 31
rect 325 50 329 55
rect 334 55 340 64
rect 375 62 377 64
rect 379 62 381 64
rect 375 61 381 62
rect 410 62 412 64
rect 414 62 416 64
rect 334 53 336 55
rect 338 53 340 55
rect 410 57 416 62
rect 432 62 434 64
rect 436 62 438 64
rect 410 55 412 57
rect 414 55 416 57
rect 410 54 416 55
rect 423 56 427 58
rect 423 54 424 56
rect 426 54 427 56
rect 432 57 438 62
rect 432 55 434 57
rect 436 55 438 57
rect 432 54 438 55
rect 464 62 466 64
rect 468 62 470 64
rect 464 57 470 62
rect 486 62 488 64
rect 490 62 492 64
rect 464 55 466 57
rect 468 55 470 57
rect 464 54 470 55
rect 475 56 479 58
rect 475 54 476 56
rect 478 54 479 56
rect 486 57 492 62
rect 521 62 523 64
rect 525 62 527 64
rect 521 61 527 62
rect 562 62 564 64
rect 566 62 568 64
rect 562 61 568 62
rect 486 55 488 57
rect 490 55 492 57
rect 486 54 492 55
rect 543 57 560 58
rect 543 55 545 57
rect 547 55 560 57
rect 543 54 560 55
rect 591 57 597 64
rect 591 55 593 57
rect 595 55 597 57
rect 591 54 597 55
rect 602 57 606 59
rect 602 55 603 57
rect 605 55 606 57
rect 334 52 340 53
rect 325 48 326 50
rect 328 49 329 50
rect 328 48 342 49
rect 325 45 342 48
rect 276 24 294 25
rect 276 22 278 24
rect 280 22 294 24
rect 276 21 294 22
rect 338 33 342 45
rect 338 31 339 33
rect 341 31 342 33
rect 338 26 342 31
rect 330 22 342 26
rect 330 18 334 22
rect 345 19 346 21
rect 216 15 217 17
rect 219 16 241 17
rect 219 15 237 16
rect 216 14 237 15
rect 239 14 241 16
rect 107 13 132 14
rect 216 13 241 14
rect 246 13 250 15
rect 314 17 334 18
rect 314 15 316 17
rect 318 15 334 17
rect 314 14 334 15
rect 380 50 404 54
rect 423 50 427 54
rect 378 46 384 50
rect 400 49 440 50
rect 400 47 424 49
rect 426 47 440 49
rect 378 36 382 46
rect 388 45 392 47
rect 400 46 440 47
rect 388 43 389 45
rect 391 43 392 45
rect 388 42 392 43
rect 378 34 379 36
rect 381 34 382 36
rect 378 32 382 34
rect 385 38 392 42
rect 385 27 389 38
rect 428 33 432 38
rect 428 31 429 33
rect 431 31 432 33
rect 371 26 389 27
rect 371 24 373 26
rect 375 25 389 26
rect 375 24 400 25
rect 371 23 396 24
rect 385 22 396 23
rect 398 22 400 24
rect 385 21 400 22
rect 405 24 409 26
rect 405 22 406 24
rect 408 22 409 24
rect 405 17 409 22
rect 428 29 432 31
rect 436 35 440 46
rect 436 33 442 35
rect 436 31 439 33
rect 441 31 442 33
rect 436 29 442 31
rect 436 26 440 29
rect 420 22 440 26
rect 420 18 424 22
rect 384 16 406 17
rect 375 13 379 15
rect 384 14 386 16
rect 388 15 406 16
rect 408 15 409 17
rect 388 14 409 15
rect 414 17 424 18
rect 414 15 416 17
rect 418 15 424 17
rect 414 14 424 15
rect 475 50 479 54
rect 498 50 522 54
rect 462 49 502 50
rect 462 47 476 49
rect 478 47 502 49
rect 462 46 502 47
rect 462 35 466 46
rect 510 45 514 47
rect 518 46 524 50
rect 510 43 511 45
rect 513 43 514 45
rect 510 42 514 43
rect 510 38 517 42
rect 460 33 466 35
rect 460 31 461 33
rect 463 31 466 33
rect 460 29 466 31
rect 470 33 474 38
rect 470 31 471 33
rect 473 31 474 33
rect 470 29 474 31
rect 462 26 466 29
rect 462 22 482 26
rect 478 18 482 22
rect 513 27 517 38
rect 520 36 524 46
rect 520 34 521 36
rect 523 34 524 36
rect 520 32 524 34
rect 513 26 531 27
rect 493 24 497 26
rect 513 25 527 26
rect 493 22 494 24
rect 496 22 497 24
rect 478 17 488 18
rect 478 15 484 17
rect 486 15 488 17
rect 478 14 488 15
rect 493 17 497 22
rect 502 24 527 25
rect 529 24 531 26
rect 502 22 504 24
rect 506 23 531 24
rect 556 50 560 54
rect 556 46 571 50
rect 546 37 552 38
rect 506 22 517 23
rect 502 21 517 22
rect 567 33 571 46
rect 574 43 575 54
rect 567 31 568 33
rect 570 31 571 33
rect 567 25 571 31
rect 602 50 606 55
rect 611 55 617 64
rect 651 62 653 64
rect 655 62 657 64
rect 651 61 657 62
rect 686 62 688 64
rect 690 62 692 64
rect 611 53 613 55
rect 615 53 617 55
rect 686 57 692 62
rect 708 62 710 64
rect 712 62 714 64
rect 686 55 688 57
rect 690 55 692 57
rect 686 54 692 55
rect 699 56 703 58
rect 699 54 700 56
rect 702 54 703 56
rect 708 57 714 62
rect 708 55 710 57
rect 712 55 714 57
rect 708 54 714 55
rect 740 62 742 64
rect 744 62 746 64
rect 740 57 746 62
rect 762 62 764 64
rect 766 62 768 64
rect 740 55 742 57
rect 744 55 746 57
rect 740 54 746 55
rect 751 56 755 58
rect 751 54 752 56
rect 754 54 755 56
rect 762 57 768 62
rect 797 62 799 64
rect 801 62 803 64
rect 797 61 803 62
rect 838 62 840 64
rect 842 62 844 64
rect 838 61 844 62
rect 762 55 764 57
rect 766 55 768 57
rect 762 54 768 55
rect 819 57 836 58
rect 819 55 821 57
rect 823 55 836 57
rect 819 54 836 55
rect 867 57 873 64
rect 867 55 869 57
rect 871 55 873 57
rect 867 54 873 55
rect 878 57 882 59
rect 878 55 879 57
rect 881 55 882 57
rect 611 52 617 53
rect 602 48 603 50
rect 605 49 606 50
rect 605 48 619 49
rect 602 45 619 48
rect 553 24 571 25
rect 553 22 555 24
rect 557 22 571 24
rect 553 21 571 22
rect 615 33 619 45
rect 615 31 616 33
rect 618 31 619 33
rect 615 26 619 31
rect 607 22 619 26
rect 607 18 611 22
rect 622 19 623 21
rect 493 15 494 17
rect 496 16 518 17
rect 496 15 514 16
rect 493 14 514 15
rect 516 14 518 16
rect 384 13 409 14
rect 493 13 518 14
rect 523 13 527 15
rect 591 17 611 18
rect 591 15 593 17
rect 595 15 611 17
rect 591 14 611 15
rect 656 50 680 54
rect 699 50 703 54
rect 654 46 660 50
rect 676 49 716 50
rect 676 47 700 49
rect 702 47 716 49
rect 654 36 658 46
rect 664 45 668 47
rect 676 46 716 47
rect 664 43 665 45
rect 667 43 668 45
rect 664 42 668 43
rect 654 34 655 36
rect 657 34 658 36
rect 654 32 658 34
rect 661 38 668 42
rect 661 27 665 38
rect 704 33 708 38
rect 704 31 705 33
rect 707 31 708 33
rect 647 26 665 27
rect 647 24 649 26
rect 651 25 665 26
rect 651 24 676 25
rect 647 23 672 24
rect 661 22 672 23
rect 674 22 676 24
rect 661 21 676 22
rect 681 24 685 26
rect 681 22 682 24
rect 684 22 685 24
rect 681 17 685 22
rect 704 29 708 31
rect 712 35 716 46
rect 712 33 718 35
rect 712 31 715 33
rect 717 31 718 33
rect 712 29 718 31
rect 712 26 716 29
rect 696 22 716 26
rect 696 18 700 22
rect 660 16 682 17
rect 651 13 655 15
rect 660 14 662 16
rect 664 15 682 16
rect 684 15 685 17
rect 664 14 685 15
rect 690 17 700 18
rect 690 15 692 17
rect 694 15 700 17
rect 690 14 700 15
rect 751 50 755 54
rect 774 50 798 54
rect 738 49 778 50
rect 738 47 752 49
rect 754 47 778 49
rect 738 46 778 47
rect 738 35 742 46
rect 786 45 790 47
rect 794 46 800 50
rect 786 43 787 45
rect 789 43 790 45
rect 786 42 790 43
rect 786 38 793 42
rect 736 33 742 35
rect 736 31 737 33
rect 739 31 742 33
rect 736 29 742 31
rect 746 33 750 38
rect 746 31 747 33
rect 749 31 750 33
rect 746 29 750 31
rect 738 26 742 29
rect 738 22 758 26
rect 754 18 758 22
rect 789 27 793 38
rect 796 36 800 46
rect 796 34 797 36
rect 799 34 800 36
rect 796 32 800 34
rect 789 26 807 27
rect 769 24 773 26
rect 789 25 803 26
rect 769 22 770 24
rect 772 22 773 24
rect 754 17 764 18
rect 754 15 760 17
rect 762 15 764 17
rect 754 14 764 15
rect 769 17 773 22
rect 778 24 803 25
rect 805 24 807 26
rect 778 22 780 24
rect 782 23 807 24
rect 832 50 836 54
rect 832 46 847 50
rect 822 37 828 38
rect 782 22 793 23
rect 778 21 793 22
rect 843 33 847 46
rect 850 43 851 54
rect 843 31 844 33
rect 846 31 847 33
rect 843 25 847 31
rect 878 50 882 55
rect 887 55 893 64
rect 928 62 930 64
rect 932 62 934 64
rect 928 61 934 62
rect 963 62 965 64
rect 967 62 969 64
rect 887 53 889 55
rect 891 53 893 55
rect 963 57 969 62
rect 985 62 987 64
rect 989 62 991 64
rect 963 55 965 57
rect 967 55 969 57
rect 963 54 969 55
rect 976 56 980 58
rect 976 54 977 56
rect 979 54 980 56
rect 985 57 991 62
rect 985 55 987 57
rect 989 55 991 57
rect 985 54 991 55
rect 1017 62 1019 64
rect 1021 62 1023 64
rect 1017 57 1023 62
rect 1039 62 1041 64
rect 1043 62 1045 64
rect 1017 55 1019 57
rect 1021 55 1023 57
rect 1017 54 1023 55
rect 1028 56 1032 58
rect 1028 54 1029 56
rect 1031 54 1032 56
rect 1039 57 1045 62
rect 1074 62 1076 64
rect 1078 62 1080 64
rect 1074 61 1080 62
rect 1115 62 1117 64
rect 1119 62 1121 64
rect 1115 61 1121 62
rect 1039 55 1041 57
rect 1043 55 1045 57
rect 1039 54 1045 55
rect 1096 57 1113 58
rect 1096 55 1098 57
rect 1100 55 1113 57
rect 1096 54 1113 55
rect 887 52 893 53
rect 878 48 879 50
rect 881 49 882 50
rect 881 48 895 49
rect 878 45 895 48
rect 829 24 847 25
rect 829 22 831 24
rect 833 22 847 24
rect 829 21 847 22
rect 891 33 895 45
rect 891 31 892 33
rect 894 31 895 33
rect 891 26 895 31
rect 883 22 895 26
rect 883 18 887 22
rect 898 19 899 21
rect 769 15 770 17
rect 772 16 794 17
rect 772 15 790 16
rect 769 14 790 15
rect 792 14 794 16
rect 660 13 685 14
rect 769 13 794 14
rect 799 13 803 15
rect 867 17 887 18
rect 867 15 869 17
rect 871 15 887 17
rect 867 14 887 15
rect 933 50 957 54
rect 976 50 980 54
rect 931 46 937 50
rect 953 49 993 50
rect 953 47 977 49
rect 979 47 993 49
rect 931 36 935 46
rect 941 45 945 47
rect 953 46 993 47
rect 941 43 942 45
rect 944 43 945 45
rect 941 42 945 43
rect 931 34 932 36
rect 934 34 935 36
rect 931 32 935 34
rect 938 38 945 42
rect 938 27 942 38
rect 981 33 985 38
rect 981 31 982 33
rect 984 31 985 33
rect 924 26 942 27
rect 924 24 926 26
rect 928 25 942 26
rect 928 24 953 25
rect 924 23 949 24
rect 938 22 949 23
rect 951 22 953 24
rect 938 21 953 22
rect 958 24 962 26
rect 958 22 959 24
rect 961 22 962 24
rect 958 17 962 22
rect 981 29 985 31
rect 989 35 993 46
rect 989 33 995 35
rect 989 31 992 33
rect 994 31 995 33
rect 989 29 995 31
rect 989 26 993 29
rect 973 22 993 26
rect 973 18 977 22
rect 937 16 959 17
rect 928 13 932 15
rect 937 14 939 16
rect 941 15 959 16
rect 961 15 962 17
rect 941 14 962 15
rect 967 17 977 18
rect 967 15 969 17
rect 971 15 977 17
rect 967 14 977 15
rect 1028 50 1032 54
rect 1051 50 1075 54
rect 1015 49 1055 50
rect 1015 47 1029 49
rect 1031 47 1055 49
rect 1015 46 1055 47
rect 1015 35 1019 46
rect 1063 45 1067 47
rect 1071 46 1077 50
rect 1063 43 1064 45
rect 1066 43 1067 45
rect 1063 42 1067 43
rect 1063 38 1070 42
rect 1013 33 1019 35
rect 1013 31 1014 33
rect 1016 31 1019 33
rect 1013 29 1019 31
rect 1023 33 1027 38
rect 1023 31 1024 33
rect 1026 31 1027 33
rect 1023 29 1027 31
rect 1015 26 1019 29
rect 1015 22 1035 26
rect 1031 18 1035 22
rect 1066 27 1070 38
rect 1073 36 1077 46
rect 1073 34 1074 36
rect 1076 34 1077 36
rect 1073 32 1077 34
rect 1066 26 1084 27
rect 1046 24 1050 26
rect 1066 25 1080 26
rect 1046 22 1047 24
rect 1049 22 1050 24
rect 1031 17 1041 18
rect 1031 15 1037 17
rect 1039 15 1041 17
rect 1031 14 1041 15
rect 1046 17 1050 22
rect 1055 24 1080 25
rect 1082 24 1084 26
rect 1055 22 1057 24
rect 1059 23 1084 24
rect 1059 22 1070 23
rect 1055 21 1070 22
rect 1109 50 1113 54
rect 1109 46 1124 50
rect 1099 37 1105 38
rect 1120 33 1124 46
rect 1127 43 1128 54
rect 1120 31 1121 33
rect 1123 31 1124 33
rect 1120 25 1124 31
rect 1106 24 1124 25
rect 1106 22 1108 24
rect 1110 22 1124 24
rect 1106 21 1124 22
rect 1046 15 1047 17
rect 1049 16 1071 17
rect 1049 15 1067 16
rect 1046 14 1067 15
rect 1069 14 1071 16
rect 937 13 962 14
rect 1046 13 1071 14
rect 1076 13 1080 15
rect -204 11 -203 13
rect -201 11 -200 13
rect -56 11 -55 13
rect -53 11 -52 13
rect -204 8 -200 11
rect -148 10 -142 11
rect -148 8 -146 10
rect -144 8 -142 10
rect -114 10 -108 11
rect -114 8 -112 10
rect -110 8 -108 10
rect -56 8 -52 11
rect -36 11 -30 12
rect -36 9 -34 11
rect -32 9 -30 11
rect -36 8 -30 9
rect -17 11 -11 12
rect -17 9 -15 11
rect -13 9 -11 11
rect -17 8 -11 9
rect 98 11 99 13
rect 101 11 102 13
rect 246 11 247 13
rect 249 11 250 13
rect 98 8 102 11
rect 154 10 160 11
rect 154 8 156 10
rect 158 8 160 10
rect 188 10 194 11
rect 188 8 190 10
rect 192 8 194 10
rect 246 8 250 11
rect 266 11 272 12
rect 266 9 268 11
rect 270 9 272 11
rect 266 8 272 9
rect 285 11 291 12
rect 285 9 287 11
rect 289 9 291 11
rect 285 8 291 9
rect 375 11 376 13
rect 378 11 379 13
rect 523 11 524 13
rect 526 11 527 13
rect 375 8 379 11
rect 431 10 437 11
rect 431 8 433 10
rect 435 8 437 10
rect 465 10 471 11
rect 465 8 467 10
rect 469 8 471 10
rect 523 8 527 11
rect 543 11 549 12
rect 543 9 545 11
rect 547 9 549 11
rect 543 8 549 9
rect 562 11 568 12
rect 562 9 564 11
rect 566 9 568 11
rect 562 8 568 9
rect 651 11 652 13
rect 654 11 655 13
rect 799 11 800 13
rect 802 11 803 13
rect 651 8 655 11
rect 707 10 713 11
rect 707 8 709 10
rect 711 8 713 10
rect 741 10 747 11
rect 741 8 743 10
rect 745 8 747 10
rect 799 8 803 11
rect 819 11 825 12
rect 819 9 821 11
rect 823 9 825 11
rect 819 8 825 9
rect 838 11 844 12
rect 838 9 840 11
rect 842 9 844 11
rect 838 8 844 9
rect 928 11 929 13
rect 931 11 932 13
rect 1076 11 1077 13
rect 1079 11 1080 13
rect 928 8 932 11
rect 984 10 990 11
rect 984 8 986 10
rect 988 8 990 10
rect 1018 10 1024 11
rect 1018 8 1020 10
rect 1022 8 1024 10
rect 1076 8 1080 11
rect 1096 11 1102 12
rect 1096 9 1098 11
rect 1100 9 1102 11
rect 1096 8 1102 9
rect 1115 11 1121 12
rect 1115 9 1117 11
rect 1119 9 1121 11
rect 1115 8 1121 9
rect -143 -16 -112 -12
rect -152 -25 -151 -19
rect -143 -20 -139 -16
rect -116 -18 -115 -16
rect -113 -18 -112 -16
rect -116 -20 -112 -18
rect -148 -24 -139 -20
rect -148 -31 -144 -24
rect -148 -33 -147 -31
rect -145 -33 -144 -31
rect -91 -16 -60 -12
rect -148 -45 -144 -33
rect -148 -47 -131 -45
rect -148 -49 -134 -47
rect -132 -49 -131 -47
rect -135 -52 -131 -49
rect -100 -25 -99 -19
rect -91 -20 -87 -16
rect -64 -18 -63 -16
rect -61 -18 -60 -16
rect -64 -20 -60 -18
rect -96 -24 -87 -20
rect -96 -31 -92 -24
rect -96 -33 -95 -31
rect -93 -33 -92 -31
rect -39 -16 -8 -12
rect -96 -45 -92 -33
rect -96 -47 -79 -45
rect -96 -49 -82 -47
rect -80 -49 -79 -47
rect -83 -52 -79 -49
rect -48 -25 -47 -19
rect -39 -20 -35 -16
rect -12 -18 -11 -16
rect -9 -18 -8 -16
rect -12 -20 -8 -18
rect -44 -24 -35 -20
rect -44 -31 -40 -24
rect -44 -33 -43 -31
rect -41 -33 -40 -31
rect 13 -16 44 -12
rect -44 -45 -40 -33
rect -44 -47 -27 -45
rect -44 -49 -30 -47
rect -28 -49 -27 -47
rect -31 -52 -27 -49
rect 4 -25 5 -19
rect 13 -20 17 -16
rect 40 -18 41 -16
rect 43 -18 44 -16
rect 40 -20 44 -18
rect 8 -24 17 -20
rect 8 -31 12 -24
rect 8 -33 9 -31
rect 11 -33 12 -31
rect 65 -16 96 -12
rect 8 -45 12 -33
rect 8 -47 25 -45
rect 8 -49 22 -47
rect 24 -49 25 -47
rect 21 -52 25 -49
rect 56 -25 57 -19
rect 65 -20 69 -16
rect 92 -18 93 -16
rect 95 -18 96 -16
rect 92 -20 96 -18
rect 60 -24 69 -20
rect 60 -31 64 -24
rect 60 -33 61 -31
rect 63 -33 64 -31
rect 118 -16 149 -12
rect 60 -45 64 -33
rect 60 -47 77 -45
rect 60 -49 74 -47
rect 76 -49 77 -47
rect 73 -52 77 -49
rect 109 -25 110 -19
rect 118 -20 122 -16
rect 145 -18 146 -16
rect 148 -18 149 -16
rect 145 -20 149 -18
rect 113 -24 122 -20
rect 113 -31 117 -24
rect 113 -33 114 -31
rect 116 -33 117 -31
rect 172 -21 178 -7
rect 172 -23 174 -21
rect 176 -23 178 -21
rect 172 -24 178 -23
rect 192 -21 198 -7
rect 192 -23 194 -21
rect 196 -23 198 -21
rect 192 -24 198 -23
rect 212 -21 218 -7
rect 212 -23 214 -21
rect 216 -23 218 -21
rect 212 -24 218 -23
rect 234 -21 240 -7
rect 234 -23 236 -21
rect 238 -23 240 -21
rect 234 -24 240 -23
rect 256 -21 262 -7
rect 256 -23 258 -21
rect 260 -23 262 -21
rect 256 -24 262 -23
rect 278 -21 284 -7
rect 278 -23 280 -21
rect 282 -23 284 -21
rect 278 -24 284 -23
rect 306 -16 337 -12
rect 113 -45 117 -33
rect 297 -25 298 -19
rect 306 -20 310 -16
rect 333 -18 334 -16
rect 336 -18 337 -16
rect 333 -20 337 -18
rect 301 -24 310 -20
rect 113 -47 130 -45
rect 113 -49 127 -47
rect 129 -49 130 -47
rect 126 -52 130 -49
rect 301 -31 305 -24
rect 301 -33 302 -31
rect 304 -33 305 -31
rect 359 -16 390 -12
rect 301 -45 305 -33
rect 301 -47 318 -45
rect 301 -49 315 -47
rect 317 -49 318 -47
rect 314 -52 318 -49
rect 350 -25 351 -19
rect 359 -20 363 -16
rect 386 -18 387 -16
rect 389 -18 390 -16
rect 386 -20 390 -18
rect 354 -24 363 -20
rect 354 -31 358 -24
rect 354 -33 355 -31
rect 357 -33 358 -31
rect 411 -16 442 -12
rect 354 -45 358 -33
rect 354 -47 371 -45
rect 354 -49 368 -47
rect 370 -49 371 -47
rect 367 -52 371 -49
rect 402 -25 403 -19
rect 411 -20 415 -16
rect 438 -18 439 -16
rect 441 -18 442 -16
rect 438 -20 442 -18
rect 406 -24 415 -20
rect 406 -31 410 -24
rect 406 -33 407 -31
rect 409 -33 410 -31
rect 463 -16 494 -12
rect 406 -45 410 -33
rect 406 -47 423 -45
rect 406 -49 420 -47
rect 422 -49 423 -47
rect 419 -52 423 -49
rect 454 -25 455 -19
rect 463 -20 467 -16
rect 490 -18 491 -16
rect 493 -18 494 -16
rect 490 -20 494 -18
rect 458 -24 467 -20
rect 458 -31 462 -24
rect 458 -33 459 -31
rect 461 -33 462 -31
rect 515 -16 546 -12
rect 458 -45 462 -33
rect 458 -47 475 -45
rect 458 -49 472 -47
rect 474 -49 475 -47
rect 471 -52 475 -49
rect 506 -25 507 -19
rect 515 -20 519 -16
rect 542 -18 543 -16
rect 545 -18 546 -16
rect 542 -20 546 -18
rect 510 -24 519 -20
rect 510 -31 514 -24
rect 510 -33 511 -31
rect 513 -33 514 -31
rect 567 -21 573 -7
rect 567 -23 569 -21
rect 571 -23 573 -21
rect 567 -24 573 -23
rect 588 -21 594 -7
rect 588 -23 590 -21
rect 592 -23 594 -21
rect 588 -24 594 -23
rect 614 -16 645 -12
rect 510 -45 514 -33
rect 510 -47 527 -45
rect 510 -49 524 -47
rect 526 -49 527 -47
rect 523 -52 527 -49
rect 605 -25 606 -19
rect 614 -20 618 -16
rect 641 -18 642 -16
rect 644 -18 645 -16
rect 641 -20 645 -18
rect 609 -24 618 -20
rect 609 -31 613 -24
rect 609 -33 610 -31
rect 612 -33 613 -31
rect 667 -16 698 -12
rect 609 -45 613 -33
rect 609 -47 626 -45
rect 609 -49 623 -47
rect 625 -49 626 -47
rect 622 -52 626 -49
rect 658 -25 659 -19
rect 667 -20 671 -16
rect 694 -18 695 -16
rect 697 -18 698 -16
rect 694 -20 698 -18
rect 662 -24 671 -20
rect 662 -31 666 -24
rect 662 -33 663 -31
rect 665 -33 666 -31
rect 719 -16 750 -12
rect 662 -45 666 -33
rect 662 -47 679 -45
rect 662 -49 676 -47
rect 678 -49 679 -47
rect 675 -52 679 -49
rect 710 -25 711 -19
rect 719 -20 723 -16
rect 746 -18 747 -16
rect 749 -18 750 -16
rect 746 -20 750 -18
rect 714 -24 723 -20
rect 714 -31 718 -24
rect 714 -33 715 -31
rect 717 -33 718 -31
rect 771 -16 802 -12
rect 714 -45 718 -33
rect 714 -47 731 -45
rect 714 -49 728 -47
rect 730 -49 731 -47
rect 727 -52 731 -49
rect 762 -25 763 -19
rect 771 -20 775 -16
rect 798 -18 799 -16
rect 801 -18 802 -16
rect 798 -20 802 -18
rect 766 -24 775 -20
rect 766 -31 770 -24
rect 766 -33 767 -31
rect 769 -33 770 -31
rect 823 -16 854 -12
rect 766 -45 770 -33
rect 766 -47 783 -45
rect 766 -49 780 -47
rect 782 -49 783 -47
rect 779 -52 783 -49
rect 814 -25 815 -19
rect 823 -20 827 -16
rect 850 -18 851 -16
rect 853 -18 854 -16
rect 850 -20 854 -18
rect 818 -24 827 -20
rect 818 -31 822 -24
rect 818 -33 819 -31
rect 821 -33 822 -31
rect 875 -16 906 -12
rect 818 -45 822 -33
rect 818 -47 835 -45
rect 818 -49 832 -47
rect 834 -49 835 -47
rect 831 -52 835 -49
rect 866 -25 867 -19
rect 875 -20 879 -16
rect 902 -18 903 -16
rect 905 -18 906 -16
rect 902 -20 906 -18
rect 870 -24 879 -20
rect 870 -31 874 -24
rect 870 -33 871 -31
rect 873 -33 874 -31
rect 928 -16 959 -12
rect 870 -45 874 -33
rect 870 -47 887 -45
rect 870 -49 884 -47
rect 886 -49 887 -47
rect 883 -52 887 -49
rect 919 -25 920 -19
rect 928 -20 932 -16
rect 955 -18 956 -16
rect 958 -18 959 -16
rect 955 -20 959 -18
rect 923 -24 932 -20
rect 923 -31 927 -24
rect 923 -33 924 -31
rect 926 -33 927 -31
rect 982 -16 1013 -12
rect 923 -45 927 -33
rect 923 -47 940 -45
rect 923 -49 937 -47
rect 939 -49 940 -47
rect 936 -52 940 -49
rect 973 -25 974 -19
rect 982 -20 986 -16
rect 1009 -18 1010 -16
rect 1012 -18 1013 -16
rect 1009 -20 1013 -18
rect 977 -24 986 -20
rect 977 -31 981 -24
rect 977 -33 978 -31
rect 980 -33 981 -31
rect 1037 -16 1068 -12
rect 977 -45 981 -33
rect 977 -47 994 -45
rect 977 -49 991 -47
rect 993 -49 994 -47
rect 990 -52 994 -49
rect 1028 -25 1029 -19
rect 1037 -20 1041 -16
rect 1064 -18 1065 -16
rect 1067 -18 1068 -16
rect 1064 -20 1068 -18
rect 1032 -24 1041 -20
rect 1032 -31 1036 -24
rect 1032 -33 1033 -31
rect 1035 -33 1036 -31
rect 1090 -16 1121 -12
rect 1032 -45 1036 -33
rect 1032 -47 1049 -45
rect 1032 -49 1046 -47
rect 1048 -49 1049 -47
rect 1045 -52 1049 -49
rect 1081 -25 1082 -19
rect 1090 -20 1094 -16
rect 1117 -18 1118 -16
rect 1120 -18 1121 -16
rect 1117 -20 1121 -18
rect 1085 -24 1094 -20
rect 1085 -31 1089 -24
rect 1085 -33 1086 -31
rect 1088 -33 1089 -31
rect 1085 -45 1089 -33
rect 1085 -47 1102 -45
rect 1085 -49 1099 -47
rect 1101 -49 1102 -47
rect 1098 -52 1102 -49
rect -135 -53 -108 -52
rect -135 -55 -112 -53
rect -110 -55 -108 -53
rect -135 -56 -108 -55
rect -83 -53 -56 -52
rect -83 -55 -60 -53
rect -58 -55 -56 -53
rect -83 -56 -56 -55
rect -31 -53 -4 -52
rect -31 -55 -8 -53
rect -6 -55 -4 -53
rect -31 -56 -4 -55
rect 21 -53 48 -52
rect 21 -55 44 -53
rect 46 -55 48 -53
rect 21 -56 48 -55
rect 73 -53 100 -52
rect 73 -55 96 -53
rect 98 -55 100 -53
rect 73 -56 100 -55
rect 126 -53 153 -52
rect 126 -55 149 -53
rect 151 -55 153 -53
rect 126 -56 153 -55
rect 314 -53 341 -52
rect 314 -55 337 -53
rect 339 -55 341 -53
rect 314 -56 341 -55
rect 367 -53 394 -52
rect 367 -55 390 -53
rect 392 -55 394 -53
rect 367 -56 394 -55
rect 419 -53 446 -52
rect 419 -55 442 -53
rect 444 -55 446 -53
rect 419 -56 446 -55
rect 471 -53 498 -52
rect 471 -55 494 -53
rect 496 -55 498 -53
rect 471 -56 498 -55
rect 523 -53 550 -52
rect 523 -55 546 -53
rect 548 -55 550 -53
rect 523 -56 550 -55
rect 622 -53 649 -52
rect 622 -55 645 -53
rect 647 -55 649 -53
rect 622 -56 649 -55
rect 675 -53 702 -52
rect 675 -55 698 -53
rect 700 -55 702 -53
rect 675 -56 702 -55
rect 727 -53 754 -52
rect 727 -55 750 -53
rect 752 -55 754 -53
rect 727 -56 754 -55
rect 779 -53 806 -52
rect 779 -55 802 -53
rect 804 -55 806 -53
rect 779 -56 806 -55
rect 831 -53 858 -52
rect 831 -55 854 -53
rect 856 -55 858 -53
rect 831 -56 858 -55
rect 883 -53 910 -52
rect 883 -55 906 -53
rect 908 -55 910 -53
rect 883 -56 910 -55
rect 936 -53 963 -52
rect 936 -55 959 -53
rect 961 -55 963 -53
rect 936 -56 963 -55
rect 990 -53 1017 -52
rect 990 -55 1013 -53
rect 1015 -55 1017 -53
rect 990 -56 1017 -55
rect 1045 -53 1072 -52
rect 1045 -55 1068 -53
rect 1070 -55 1072 -53
rect 1045 -56 1072 -55
rect 1098 -53 1125 -52
rect 1098 -55 1121 -53
rect 1123 -55 1125 -53
rect 1098 -56 1125 -55
<< via1 >>
rect 98 356 100 358
rect -276 342 -274 344
rect -265 320 -263 322
rect -226 320 -224 322
rect -274 311 -272 313
rect -265 310 -263 312
rect -182 320 -180 322
rect -157 319 -155 321
rect -214 311 -212 313
rect -133 319 -131 321
rect -123 332 -121 334
rect -104 327 -102 329
rect -92 311 -90 313
rect -35 332 -33 334
rect -35 319 -33 321
rect 8 330 10 332
rect -3 315 -1 317
rect -44 307 -42 309
rect 16 310 18 312
rect 48 336 50 338
rect 40 324 42 326
rect 56 313 58 315
rect 80 319 82 321
rect 120 327 122 329
rect 138 319 140 321
rect 88 311 90 313
rect 169 319 171 321
rect 179 332 181 334
rect 209 327 211 329
rect 210 311 212 313
rect 267 336 269 338
rect 267 319 269 321
rect 315 332 317 334
rect 299 315 301 317
rect 258 307 260 309
rect 332 319 334 321
rect 347 324 349 326
rect 397 327 399 329
rect 415 319 417 321
rect 365 311 367 313
rect 446 319 448 321
rect 456 332 458 334
rect 486 327 488 329
rect 487 311 489 313
rect 544 336 546 338
rect 544 319 546 321
rect 592 332 594 334
rect 576 315 578 317
rect 535 307 537 309
rect 609 319 611 321
rect 624 324 626 326
rect 673 327 675 329
rect 691 319 693 321
rect 641 311 643 313
rect 722 319 724 321
rect 732 332 734 334
rect 762 327 764 329
rect 763 311 765 313
rect 820 336 822 338
rect 811 308 813 310
rect 820 319 822 321
rect 868 332 870 334
rect 852 315 854 317
rect 885 319 887 321
rect 900 324 902 326
rect 950 327 952 329
rect 968 319 970 321
rect 918 311 920 313
rect 999 319 1001 321
rect 1009 332 1011 334
rect 1039 327 1041 329
rect 1040 311 1042 313
rect 1097 336 1099 338
rect 1097 319 1099 321
rect 1129 315 1131 317
rect 1088 306 1090 308
rect 211 290 213 292
rect 488 290 490 292
rect 764 290 766 292
rect 1041 290 1043 292
rect 164 288 166 290
rect -265 264 -263 266
rect -226 254 -224 256
rect -281 237 -279 239
rect -214 263 -212 265
rect -182 254 -180 256
rect -164 255 -162 257
rect -133 255 -131 257
rect -92 263 -90 265
rect -123 242 -121 244
rect -44 263 -42 265
rect -88 247 -86 249
rect -35 255 -33 257
rect -35 242 -33 244
rect 16 259 18 261
rect -3 247 -1 249
rect 16 247 18 249
rect 56 264 58 266
rect 40 247 42 249
rect 80 255 82 257
rect 48 239 50 241
rect 88 263 90 265
rect 138 255 140 257
rect 169 255 171 257
rect 133 247 135 249
rect 210 263 212 265
rect 179 242 181 244
rect 260 269 262 271
rect 227 250 229 252
rect 267 261 269 263
rect 267 242 269 244
rect 332 255 334 257
rect 315 247 317 249
rect 347 254 349 256
rect 291 231 293 233
rect 365 263 367 265
rect 415 255 417 257
rect 446 255 448 257
rect 410 247 412 249
rect 487 263 489 265
rect 456 242 458 244
rect 537 269 539 271
rect 504 250 506 252
rect 544 261 546 263
rect 544 242 546 244
rect 609 255 611 257
rect 592 247 594 249
rect 624 254 626 256
rect 568 231 570 233
rect 641 263 643 265
rect 691 255 693 257
rect 722 255 724 257
rect 686 247 688 249
rect 763 263 765 265
rect 732 242 734 244
rect 813 269 815 271
rect 780 250 782 252
rect 820 261 822 263
rect 820 242 822 244
rect 885 255 887 257
rect 868 247 870 249
rect 900 254 902 256
rect 844 231 846 233
rect 918 263 920 265
rect 968 255 970 257
rect 999 255 1001 257
rect 963 247 965 249
rect 1090 272 1092 274
rect 1040 263 1042 265
rect 1009 242 1011 244
rect 1057 250 1059 252
rect 1097 261 1099 263
rect 1097 242 1099 244
rect 1121 231 1123 233
rect 100 216 102 218
rect -281 186 -279 188
rect -265 175 -263 177
rect -226 176 -224 178
rect -182 176 -180 178
rect -163 175 -161 177
rect -214 167 -212 169
rect -133 175 -131 177
rect -123 188 -121 190
rect -86 183 -84 185
rect -92 167 -90 169
rect -35 188 -33 190
rect -44 165 -42 167
rect -35 175 -33 177
rect 8 186 10 188
rect -3 171 -1 173
rect 40 183 42 185
rect 48 192 50 194
rect 16 167 18 169
rect 56 170 58 172
rect 80 175 82 177
rect 137 183 139 185
rect 139 175 141 177
rect 88 167 90 169
rect 169 175 171 177
rect 179 188 181 190
rect 227 183 229 185
rect 210 167 212 169
rect 267 192 269 194
rect 267 175 269 177
rect 315 187 317 189
rect 299 171 301 173
rect 332 175 334 177
rect 347 180 349 182
rect 260 159 262 161
rect 414 183 416 185
rect 416 175 418 177
rect 365 167 367 169
rect 446 175 448 177
rect 456 188 458 190
rect 504 183 506 185
rect 487 167 489 169
rect 544 192 546 194
rect 544 175 546 177
rect 592 187 594 189
rect 576 171 578 173
rect 609 175 611 177
rect 624 180 626 182
rect 537 159 539 161
rect 690 183 692 185
rect 692 175 694 177
rect 641 167 643 169
rect 722 175 724 177
rect 732 188 734 190
rect 780 183 782 185
rect 763 167 765 169
rect 820 192 822 194
rect 820 175 822 177
rect 868 187 870 189
rect 852 171 854 173
rect 885 175 887 177
rect 900 180 902 182
rect 813 159 815 161
rect 967 183 969 185
rect 969 175 971 177
rect 918 167 920 169
rect 999 175 1001 177
rect 1009 188 1011 190
rect 1057 183 1059 185
rect 1040 167 1042 169
rect 1097 192 1099 194
rect 1097 175 1099 177
rect 1129 171 1131 173
rect 1088 162 1090 164
rect 165 144 167 146
rect -265 120 -263 122
rect -226 110 -224 112
rect -281 90 -279 92
rect -214 119 -212 121
rect -182 110 -180 112
rect -157 111 -155 113
rect -133 111 -131 113
rect -92 119 -90 121
rect -123 98 -121 100
rect -44 124 -42 126
rect -88 103 -86 105
rect -35 111 -33 113
rect -35 98 -33 100
rect 16 115 18 117
rect -3 103 -1 105
rect 17 103 19 105
rect 56 119 58 121
rect 40 103 42 105
rect 80 111 82 113
rect 48 95 50 97
rect 88 119 90 121
rect 138 111 140 113
rect 169 111 171 113
rect 131 103 133 105
rect 210 119 212 121
rect 179 98 181 100
rect 260 125 262 127
rect 227 106 229 108
rect 267 117 269 119
rect 267 98 269 100
rect 332 111 334 113
rect 315 103 317 105
rect 347 107 349 109
rect 290 87 292 89
rect 365 119 367 121
rect 415 111 417 113
rect 446 111 448 113
rect 408 103 410 105
rect 487 119 489 121
rect 456 98 458 100
rect 537 125 539 127
rect 504 106 506 108
rect 544 117 546 119
rect 544 98 546 100
rect 609 111 611 113
rect 592 103 594 105
rect 624 107 626 109
rect 567 87 569 89
rect 641 119 643 121
rect 691 111 693 113
rect 722 111 724 113
rect 684 103 686 105
rect 763 119 765 121
rect 732 98 734 100
rect 813 125 815 127
rect 780 106 782 108
rect 820 117 822 119
rect 820 98 822 100
rect 885 111 887 113
rect 868 103 870 105
rect 900 107 902 109
rect 843 87 845 89
rect 918 119 920 121
rect 968 111 970 113
rect 999 111 1001 113
rect 961 103 963 105
rect 1090 127 1092 129
rect 1040 119 1042 121
rect 1009 98 1011 100
rect 1057 106 1059 108
rect 1097 117 1099 119
rect 1097 98 1099 100
rect 1120 87 1122 89
rect 99 71 101 73
rect 1069 72 1071 74
rect -282 51 -280 53
rect -265 31 -263 33
rect -226 32 -224 34
rect -182 32 -180 34
rect -163 31 -161 33
rect -214 23 -212 25
rect -133 31 -131 33
rect -123 44 -121 46
rect -88 39 -86 41
rect -92 23 -90 25
rect -35 44 -33 46
rect -44 20 -42 22
rect -35 31 -33 33
rect 8 42 10 44
rect -3 29 -1 31
rect 15 22 17 24
rect 48 48 50 50
rect 56 25 58 27
rect 80 31 82 33
rect 32 15 34 17
rect 133 39 135 41
rect 138 31 140 33
rect 88 23 90 25
rect 169 31 171 33
rect 179 44 181 46
rect 226 39 228 41
rect 210 23 212 25
rect 267 48 269 50
rect 258 21 260 23
rect 267 31 269 33
rect 315 47 317 49
rect 299 31 301 33
rect 332 31 334 33
rect 347 37 349 39
rect 410 39 412 41
rect 415 31 417 33
rect 365 23 367 25
rect 446 31 448 33
rect 456 44 458 46
rect 503 39 505 41
rect 487 23 489 25
rect 544 48 546 50
rect 535 21 537 23
rect 544 31 546 33
rect 592 47 594 49
rect 576 31 578 33
rect 609 31 611 33
rect 624 37 626 39
rect 686 39 688 41
rect 691 31 693 33
rect 641 23 643 25
rect 722 31 724 33
rect 732 44 734 46
rect 779 39 781 41
rect 763 23 765 25
rect 820 48 822 50
rect 811 21 813 23
rect 820 31 822 33
rect 868 47 870 49
rect 852 31 854 33
rect 885 31 887 33
rect 900 37 902 39
rect 963 39 965 41
rect 968 31 970 33
rect 918 23 920 25
rect 999 31 1001 33
rect 1009 44 1011 46
rect 1056 39 1058 41
rect 1040 23 1042 25
rect 1097 48 1099 50
rect 1097 31 1099 33
rect 1129 28 1131 30
rect 1088 18 1090 20
rect 134 2 136 4
rect 164 3 166 5
rect -131 -23 -129 -21
rect -114 -40 -112 -38
rect -120 -48 -118 -46
rect -79 -23 -77 -21
rect -62 -40 -60 -38
rect -69 -48 -67 -46
rect -27 -23 -25 -21
rect -10 -40 -8 -38
rect -16 -48 -14 -46
rect 25 -31 27 -29
rect 42 -40 44 -38
rect 35 -48 37 -46
rect 77 -29 79 -27
rect 94 -40 96 -38
rect 87 -48 89 -46
rect 130 -24 132 -22
rect 184 -26 186 -24
rect 210 -33 212 -31
rect 230 -33 232 -31
rect 250 -33 252 -31
rect 147 -40 149 -38
rect 171 -40 173 -38
rect 277 -41 279 -39
rect 318 -24 320 -22
rect 294 -42 296 -40
rect 140 -48 142 -46
rect 163 -47 165 -45
rect 183 -47 185 -45
rect 203 -49 205 -47
rect 225 -48 227 -46
rect 247 -50 249 -48
rect 269 -51 271 -49
rect 335 -40 337 -38
rect 329 -48 331 -46
rect 368 -32 370 -30
rect 388 -40 390 -38
rect 382 -48 384 -46
rect 423 -29 425 -27
rect 440 -40 442 -38
rect 433 -48 435 -46
rect 473 -32 475 -30
rect 492 -40 494 -38
rect 486 -48 488 -46
rect 527 -28 529 -26
rect 544 -40 546 -38
rect 566 -38 568 -36
rect 587 -40 589 -38
rect 537 -48 539 -46
rect 626 -25 628 -23
rect 643 -40 645 -38
rect 643 -48 645 -46
rect 679 -23 681 -21
rect 696 -40 698 -38
rect 690 -48 692 -46
rect 731 -24 733 -22
rect 748 -40 750 -38
rect 741 -48 743 -46
rect 783 -24 785 -22
rect 800 -40 802 -38
rect 794 -48 796 -46
rect 835 -24 837 -22
rect 852 -40 854 -38
rect 845 -48 847 -46
rect 887 -24 889 -22
rect 904 -40 906 -38
rect 897 -48 899 -46
rect 940 -24 942 -22
rect 957 -40 959 -38
rect 950 -48 952 -46
rect 994 -24 996 -22
rect 1011 -40 1013 -38
rect 1002 -48 1004 -46
rect 1049 -24 1051 -22
rect 1066 -40 1068 -38
rect 1059 -48 1061 -46
rect 1102 -24 1104 -22
rect 1119 -40 1121 -38
rect 1111 -48 1113 -46
rect -151 -56 -149 -54
rect -99 -56 -97 -54
rect -47 -56 -45 -54
rect 5 -56 7 -54
rect 57 -57 59 -55
rect 110 -57 112 -55
rect 351 -57 353 -55
rect 403 -57 405 -55
rect 455 -57 457 -55
rect 507 -57 509 -55
rect 558 -54 560 -52
rect 580 -56 582 -54
rect 607 -57 609 -55
rect 659 -56 661 -54
rect 711 -57 713 -55
rect 763 -57 765 -55
rect 816 -57 818 -55
rect 867 -57 869 -55
rect 920 -57 922 -55
rect 974 -57 976 -55
rect 1030 -57 1032 -55
rect 1086 -57 1088 -55
rect 1078 -67 1080 -65
<< via2 >>
rect 90 356 92 358
rect -276 346 -274 348
rect 45 348 47 350
rect 185 348 187 350
rect 2 330 4 332
rect -131 328 -129 330
rect -112 327 -110 329
rect 215 327 217 329
rect 492 327 494 329
rect 768 327 770 329
rect 1045 327 1047 329
rect -164 319 -162 321
rect -44 311 -42 313
rect -84 287 -82 289
rect 44 313 46 315
rect 303 315 305 317
rect 262 307 264 309
rect 169 288 171 290
rect 215 290 217 292
rect 264 290 266 292
rect 323 290 325 292
rect -161 278 -159 280
rect 211 277 213 279
rect 314 277 316 279
rect -281 243 -279 245
rect -281 178 -279 180
rect -68 264 -66 266
rect 264 269 266 271
rect 2 259 4 261
rect -161 255 -159 257
rect 303 250 305 252
rect -84 247 -82 249
rect -90 216 -88 218
rect 580 315 582 317
rect 535 303 537 305
rect 343 290 345 292
rect 492 290 494 292
rect 541 290 543 292
rect 600 290 602 292
rect 348 277 350 279
rect 591 277 593 279
rect 541 269 543 271
rect 44 239 46 241
rect 89 215 91 217
rect -163 205 -161 207
rect 236 204 238 206
rect 264 204 266 206
rect 2 186 4 188
rect 323 214 325 216
rect -90 183 -88 185
rect 307 204 309 206
rect -28 165 -26 167
rect 44 170 46 172
rect 303 171 305 173
rect 580 250 582 252
rect 856 315 858 317
rect 791 308 793 310
rect 620 290 622 292
rect 768 290 770 292
rect 817 290 819 292
rect 876 290 878 292
rect 625 277 627 279
rect 817 269 819 271
rect 341 214 343 216
rect 347 205 349 207
rect 541 204 543 206
rect 600 214 602 216
rect 584 204 586 206
rect -84 143 -82 145
rect 332 165 334 167
rect 169 143 171 145
rect 264 142 266 144
rect 324 142 326 144
rect -164 132 -162 134
rect 253 133 255 135
rect 311 133 313 135
rect -40 125 -38 127
rect -281 87 -279 89
rect -282 48 -280 50
rect 264 125 266 127
rect 2 115 4 117
rect -164 111 -162 113
rect 303 106 305 108
rect -84 103 -82 105
rect -84 70 -82 72
rect 580 171 582 173
rect 856 250 858 252
rect 1133 315 1135 317
rect 1088 297 1090 299
rect 896 290 898 292
rect 1045 290 1047 292
rect 1084 272 1086 274
rect 618 214 620 216
rect 624 205 626 207
rect 817 204 819 206
rect 876 214 878 216
rect 860 204 862 206
rect 340 142 342 144
rect 541 142 543 144
rect 601 142 603 144
rect 347 133 349 135
rect 588 133 590 135
rect 541 125 543 127
rect 44 95 46 97
rect 89 71 91 73
rect -163 60 -161 62
rect 261 61 263 63
rect 2 42 4 44
rect 323 70 325 72
rect 307 61 309 63
rect -84 39 -82 41
rect 129 39 131 41
rect 193 31 195 33
rect 303 31 305 33
rect 580 106 582 108
rect 856 171 858 173
rect 1133 250 1135 252
rect 894 214 896 216
rect 617 142 619 144
rect 817 142 819 144
rect 877 142 879 144
rect 624 133 626 135
rect 864 133 866 135
rect 817 125 819 127
rect 340 70 342 72
rect 345 62 347 64
rect 538 61 540 63
rect 856 106 858 108
rect 1133 171 1135 173
rect 893 142 895 144
rect 940 143 942 145
rect 1084 127 1086 129
rect 609 86 611 88
rect 600 70 602 72
rect 584 61 586 63
rect -13 20 -11 22
rect -131 -4 -129 -2
rect -68 -2 -66 0
rect 44 25 46 27
rect 19 22 21 24
rect 357 31 359 33
rect 580 31 582 33
rect 617 70 619 72
rect 622 62 624 64
rect 814 61 816 63
rect 876 70 878 72
rect 860 61 862 63
rect 35 16 37 18
rect 634 31 636 33
rect 856 31 858 33
rect 1133 106 1135 108
rect 893 70 895 72
rect 1074 70 1076 72
rect 885 44 887 46
rect 910 31 912 33
rect 129 2 131 4
rect 169 3 171 5
rect 672 2 674 4
rect -27 -17 -25 -15
rect 25 -25 27 -23
rect 77 -24 79 -22
rect 626 -17 628 -15
rect 791 0 793 2
rect 725 -6 727 -4
rect 887 -5 889 -3
rect 841 -18 843 -16
rect 1019 -6 1021 -4
rect 940 -19 942 -17
rect 205 -33 207 -31
rect 233 -33 235 -31
rect 299 -33 301 -31
rect 362 -32 364 -30
rect 421 -32 423 -30
rect 466 -32 468 -30
rect 527 -32 529 -30
rect 335 -37 337 -35
rect 284 -41 286 -39
rect 298 -42 300 -40
rect 171 -45 173 -43
rect 188 -47 190 -45
rect 203 -45 205 -43
rect 234 -49 236 -47
rect 247 -47 249 -45
rect 269 -48 271 -46
rect 163 -53 165 -51
rect 558 -51 560 -49
rect 1074 -67 1076 -65
<< via3 >>
rect 85 355 87 357
rect 31 348 33 350
rect 188 348 190 350
rect -164 337 -162 339
rect -51 314 -49 316
rect -281 271 -279 273
rect -60 271 -58 273
rect -6 271 -4 273
rect -281 173 -279 175
rect -277 87 -275 89
rect -282 44 -280 46
rect -24 165 -22 167
rect -40 121 -38 123
rect 265 307 267 309
rect 174 289 176 291
rect 44 271 46 273
rect 85 215 87 217
rect 173 143 175 145
rect 85 71 87 73
rect -102 -4 -100 -2
rect 24 22 26 24
rect 39 16 41 18
rect 160 31 162 33
rect 197 30 199 32
rect 174 3 176 5
rect 535 300 537 302
rect 411 288 413 290
rect 211 2 213 4
rect 237 0 239 2
rect 329 165 331 167
rect 726 286 728 288
rect 603 87 605 89
rect 550 70 552 72
rect 672 71 674 73
rect 270 61 272 63
rect 253 1 255 3
rect -23 -17 -21 -15
rect 25 -19 27 -17
rect 188 -4 190 -2
rect 163 -61 165 -59
rect 1088 287 1090 289
rect 876 44 878 46
rect 842 1 844 3
rect 517 -12 519 -10
rect 347 -24 349 -22
rect 327 -33 329 -31
rect 371 -24 373 -22
rect 458 -33 460 -31
rect 626 -9 628 -7
rect 271 -41 273 -39
rect 211 -45 213 -43
rect 238 -48 240 -46
rect 253 -47 255 -45
rect 289 -41 291 -39
rect 301 -42 303 -40
rect 335 -43 337 -41
rect 285 -54 287 -52
rect 335 -64 337 -62
<< via4 >>
rect -281 165 -279 167
rect -274 87 -272 89
rect -274 44 -272 46
rect 17 271 19 273
rect 38 271 40 273
rect -40 -1 -38 1
rect 325 164 327 166
rect 598 87 600 89
rect 870 44 872 46
rect 25 -14 27 -12
<< labels >>
rlabel alu1 108 355 108 355 1 Vdd
rlabel alu1 -280 190 -280 190 1 b2
rlabel alu1 -281 96 -281 96 1 b3
rlabel alu1 -281 46 -281 46 1 b4
rlabel alu1 53 288 53 288 1 Gnd
rlabel alu2 -157 -48 -157 -48 1 x0
rlabel alu2 -157 -40 -157 -40 1 x1
rlabel alu2 -288 312 -288 312 3 cin
rlabel alu1 -289 339 -289 339 3 b0
rlabel alu3 -289 319 -289 319 3 a0
rlabel alu3 -286 281 -286 281 3 a1
rlabel alu1 -286 231 -286 231 3 b1
rlabel alu3 -282 206 -282 206 1 a2
rlabel alu3 -284 134 -284 134 1 a3
rlabel alu3 -286 61 -286 61 3 a4
rlabel alu2 -150 -79 -150 -79 1 s0
rlabel alu2 -99 -80 -99 -80 1 s1
rlabel alu2 -47 -78 -47 -78 1 s2
rlabel alu2 5 -78 5 -78 1 s3
rlabel alu2 57 -79 57 -79 1 s4
rlabel alu2 111 -80 111 -80 1 cout
rlabel alu4 302 -77 302 -77 1 i0
rlabel alu2 352 -79 352 -79 1 i1
rlabel alu2 404 -78 404 -78 1 i2
rlabel alu2 455 -78 455 -78 1 i3
rlabel alu2 508 -78 508 -78 1 i4
rlabel alu2 608 -78 608 -78 1 p0
rlabel alu2 660 -77 660 -77 1 p1
rlabel alu2 711 -80 711 -80 1 p2
rlabel alu2 764 -78 764 -78 1 p3
rlabel alu2 817 -79 817 -79 1 p4
rlabel alu2 867 -81 867 -81 1 p5
rlabel alu2 921 -79 921 -79 1 p6
rlabel alu2 975 -78 975 -78 1 p7
rlabel alu2 1030 -78 1030 -78 1 p8
rlabel alu2 1086 -80 1086 -80 1 p9
<< end >>
